<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-1540.15,-3163.5,-316.15,-3768.5</PageViewport>
<gate>
<ID>2307</ID>
<type>AA_AND2</type>
<position>-1151,-3266</position>
<input>
<ID>IN_0</ID>2521 </input>
<input>
<ID>IN_1</ID>2526 </input>
<output>
<ID>OUT</ID>2522 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2308</ID>
<type>AA_AND2</type>
<position>-1133.5,-3267</position>
<input>
<ID>IN_0</ID>2522 </input>
<input>
<ID>IN_1</ID>2528 </input>
<output>
<ID>OUT</ID>2523 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2309</ID>
<type>AA_AND2</type>
<position>-1279.5,-3193</position>
<input>
<ID>IN_0</ID>2504 </input>
<input>
<ID>IN_1</ID>2510 </input>
<output>
<ID>OUT</ID>2505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2310</ID>
<type>BA_NAND4</type>
<position>-1111.5,-3264</position>
<input>
<ID>IN_0</ID>2527 </input>
<input>
<ID>IN_1</ID>2526 </input>
<input>
<ID>IN_2</ID>2528 </input>
<input>
<ID>IN_3</ID>2529 </input>
<output>
<ID>OUT</ID>2208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2311</ID>
<type>AE_DFF_LOW</type>
<position>-1194.5,-3309.5</position>
<input>
<ID>IN_0</ID>2524 </input>
<output>
<ID>OUT_0</ID>2530 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2312</ID>
<type>AA_AND2</type>
<position>-1262,-3194</position>
<input>
<ID>IN_0</ID>2505 </input>
<input>
<ID>IN_1</ID>2512 </input>
<output>
<ID>OUT</ID>2506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2313</ID>
<type>AE_DFF_LOW</type>
<position>-1178,-3309.5</position>
<input>
<ID>IN_0</ID>2525 </input>
<output>
<ID>OUT_0</ID>2531 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2314</ID>
<type>AE_DFF_LOW</type>
<position>-1163.5,-3309.5</position>
<input>
<ID>IN_0</ID>2527 </input>
<output>
<ID>OUT_0</ID>2532 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2315</ID>
<type>BA_NAND4</type>
<position>-1240,-3191</position>
<input>
<ID>IN_0</ID>2511 </input>
<input>
<ID>IN_1</ID>2510 </input>
<input>
<ID>IN_2</ID>2512 </input>
<input>
<ID>IN_3</ID>2513 </input>
<output>
<ID>OUT</ID>2495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2316</ID>
<type>AE_DFF_LOW</type>
<position>-1146.5,-3309.5</position>
<input>
<ID>IN_0</ID>2526 </input>
<output>
<ID>OUT_0</ID>2533 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2317</ID>
<type>AE_DFF_LOW</type>
<position>-1130.5,-3309.5</position>
<input>
<ID>IN_0</ID>2528 </input>
<output>
<ID>OUT_0</ID>2534 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2318</ID>
<type>AE_DFF_LOW</type>
<position>-1112.5,-3309.5</position>
<input>
<ID>IN_0</ID>2529 </input>
<output>
<ID>OUT_0</ID>2535 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2319</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-1092.5,-3319</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2531 </input>
<input>
<ID>IN_2</ID>2532 </input>
<input>
<ID>IN_3</ID>2533 </input>
<input>
<ID>IN_4</ID>2534 </input>
<input>
<ID>IN_5</ID>2535 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2320</ID>
<type>AA_INVERTER</type>
<position>-1205,-3216.5</position>
<input>
<ID>IN_0</ID>2494 </input>
<output>
<ID>OUT_0</ID>2537 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2321</ID>
<type>AE_DFF_LOW</type>
<position>-1323,-3236.5</position>
<input>
<ID>IN_0</ID>2507 </input>
<output>
<ID>OUT_0</ID>2514 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2322</ID>
<type>AE_DFF_LOW</type>
<position>-1306.5,-3236.5</position>
<input>
<ID>IN_0</ID>2509 </input>
<output>
<ID>OUT_0</ID>2515 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2323</ID>
<type>AE_DFF_LOW</type>
<position>-1292,-3236.5</position>
<input>
<ID>IN_0</ID>2511 </input>
<output>
<ID>OUT_0</ID>2516 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2324</ID>
<type>AE_DFF_LOW</type>
<position>-1275,-3236.5</position>
<input>
<ID>IN_0</ID>2510 </input>
<output>
<ID>OUT_0</ID>2517 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2325</ID>
<type>AE_DFF_LOW</type>
<position>-1259,-3236.5</position>
<input>
<ID>IN_0</ID>2512 </input>
<output>
<ID>OUT_0</ID>2518 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2326</ID>
<type>AE_DFF_LOW</type>
<position>-1241,-3236.5</position>
<input>
<ID>IN_0</ID>2513 </input>
<output>
<ID>OUT_0</ID>2519 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2327</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-1221,-3246</position>
<input>
<ID>IN_0</ID>2514 </input>
<input>
<ID>IN_1</ID>2515 </input>
<input>
<ID>IN_2</ID>2516 </input>
<input>
<ID>IN_3</ID>2517 </input>
<input>
<ID>IN_4</ID>2518 </input>
<input>
<ID>IN_5</ID>2519 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2328</ID>
<type>AA_AND2</type>
<position>-1358.5,-3205.5</position>
<input>
<ID>IN_0</ID>2666 </input>
<input>
<ID>IN_1</ID>2424 </input>
<output>
<ID>OUT</ID>2536 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2329</ID>
<type>AE_DFF_LOW</type>
<position>-1414.5,-3372.5</position>
<input>
<ID>IN_0</ID>2419 </input>
<output>
<ID>OUTINV_0</ID>2425 </output>
<output>
<ID>OUT_0</ID>2423 </output>
<input>
<ID>clock</ID>2421 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2330</ID>
<type>AA_TOGGLE</type>
<position>-1427,-3370.5</position>
<output>
<ID>OUT_0</ID>2419 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2331</ID>
<type>AI_XOR2</type>
<position>-870,-3592.5</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2553 </input>
<output>
<ID>OUT</ID>2396 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2332</ID>
<type>AI_XOR2</type>
<position>-856.5,-3592.5</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2555 </input>
<output>
<ID>OUT</ID>2397 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2333</ID>
<type>AA_AND2</type>
<position>-1398,-3361.5</position>
<input>
<ID>IN_0</ID>2423 </input>
<input>
<ID>IN_1</ID>2422 </input>
<output>
<ID>OUT</ID>2424 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2334</ID>
<type>AI_XOR2</type>
<position>-843.5,-3592.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2557 </input>
<output>
<ID>OUT</ID>2398 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2335</ID>
<type>AA_LABEL</type>
<position>-1431,-3361</position>
<gparam>LABEL_TEXT On/Off Switch</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2336</ID>
<type>AI_XOR2</type>
<position>-830.5,-3592.5</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2559 </input>
<output>
<ID>OUT</ID>2399 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2337</ID>
<type>AI_XOR2</type>
<position>-818,-3593</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2561 </input>
<output>
<ID>OUT</ID>2400 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2338</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1404,-3373.5</position>
<input>
<ID>IN_0</ID>2425 </input>
<output>
<ID>OUT_0</ID>2426 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2339</ID>
<type>AI_XOR2</type>
<position>-805.5,-3593</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2563 </input>
<output>
<ID>OUT</ID>2401 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2340</ID>
<type>AA_LABEL</type>
<position>-1276,-3383</position>
<gparam>LABEL_TEXT Default Power</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2341</ID>
<type>AE_DFF_LOW</type>
<position>-1364.5,-3374.5</position>
<input>
<ID>IN_0</ID>2420 </input>
<output>
<ID>OUTINV_0</ID>2422 </output>
<output>
<ID>OUT_0</ID>2478 </output>
<input>
<ID>clear</ID>2426 </input>
<input>
<ID>clock</ID>2421 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2342</ID>
<type>BB_CLOCK</type>
<position>-1379.5,-3378</position>
<output>
<ID>CLK</ID>2421 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>2343</ID>
<type>AA_AND2</type>
<position>-783,-4514.5</position>
<input>
<ID>IN_0</ID>2542 </input>
<input>
<ID>IN_1</ID>2541 </input>
<output>
<ID>OUT</ID>2545 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2344</ID>
<type>AA_TOGGLE</type>
<position>-990,-3643.5</position>
<output>
<ID>OUT_0</ID>2691 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2345</ID>
<type>AA_AND2</type>
<position>-805.5,-4537.5</position>
<input>
<ID>IN_0</ID>2545 </input>
<input>
<ID>IN_1</ID>2543 </input>
<output>
<ID>OUT</ID>2306 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2346</ID>
<type>AA_AND2</type>
<position>-959,-3710</position>
<input>
<ID>IN_0</ID>2544 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2347</ID>
<type>AA_AND2</type>
<position>-959.5,-3701.5</position>
<input>
<ID>IN_0</ID>2544 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2348</ID>
<type>AA_AND2</type>
<position>-960,-3693</position>
<input>
<ID>IN_0</ID>2544 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2643 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2349</ID>
<type>AA_AND2</type>
<position>-960.5,-3685</position>
<input>
<ID>IN_0</ID>2544 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2350</ID>
<type>AA_AND2</type>
<position>-961,-3676.5</position>
<input>
<ID>IN_0</ID>2544 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2647 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2351</ID>
<type>AA_AND2</type>
<position>-961,-3668</position>
<input>
<ID>IN_0</ID>2544 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2352</ID>
<type>AI_XOR2</type>
<position>-848.5,-4482.5</position>
<input>
<ID>IN_0</ID>2278 </input>
<input>
<ID>IN_1</ID>2547 </input>
<output>
<ID>OUT</ID>2388 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2353</ID>
<type>AA_LABEL</type>
<position>-997,-3483.5</position>
<gparam>LABEL_TEXT Zone 1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2354</ID>
<type>AI_XOR2</type>
<position>-835,-4482.5</position>
<input>
<ID>IN_0</ID>2299 </input>
<input>
<ID>IN_1</ID>2549 </input>
<output>
<ID>OUT</ID>2389 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2355</ID>
<type>AA_LABEL</type>
<position>-989.5,-3633</position>
<gparam>LABEL_TEXT Zone 2</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2356</ID>
<type>AI_XOR2</type>
<position>-822,-4482.5</position>
<input>
<ID>IN_0</ID>2300 </input>
<input>
<ID>IN_1</ID>2551 </input>
<output>
<ID>OUT</ID>2390 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2357</ID>
<type>AI_XOR2</type>
<position>-809,-4482.5</position>
<input>
<ID>IN_0</ID>2301 </input>
<input>
<ID>IN_1</ID>2566 </input>
<output>
<ID>OUT</ID>2391 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2358</ID>
<type>AI_XOR2</type>
<position>-796.5,-4483</position>
<input>
<ID>IN_0</ID>2302 </input>
<input>
<ID>IN_1</ID>2568 </input>
<output>
<ID>OUT</ID>2392 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2359</ID>
<type>AI_XOR2</type>
<position>-784,-4483</position>
<input>
<ID>IN_0</ID>2304 </input>
<input>
<ID>IN_1</ID>2570 </input>
<output>
<ID>OUT</ID>2394 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2360</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-891,-3555.5</position>
<input>
<ID>J</ID>2552 </input>
<output>
<ID>Q</ID>2553 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2652 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2361</ID>
<type>AI_XOR2</type>
<position>-757.5,-4993</position>
<input>
<ID>IN_0</ID>2326 </input>
<input>
<ID>IN_1</ID>2328 </input>
<output>
<ID>OUT</ID>2329 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2362</ID>
<type>AA_LABEL</type>
<position>-981.5,-4353</position>
<gparam>LABEL_TEXT Zone 6</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2363</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-904,-3545.5</position>
<input>
<ID>J</ID>2554 </input>
<output>
<ID>Q</ID>2555 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2652 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2364</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-917,-3534.5</position>
<input>
<ID>J</ID>2556 </input>
<output>
<ID>Q</ID>2557 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2652 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2365</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-924.5,-3525.5</position>
<input>
<ID>J</ID>2558 </input>
<output>
<ID>Q</ID>2559 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2652 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2366</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-933,-3518</position>
<input>
<ID>J</ID>2560 </input>
<output>
<ID>Q</ID>2561 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2652 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2367</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-942,-3510.5</position>
<input>
<ID>J</ID>2562 </input>
<output>
<ID>Q</ID>2563 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2652 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2368</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-901,-3712</position>
<input>
<ID>J</ID>2564 </input>
<output>
<ID>Q</ID>2640 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2651 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2369</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-799,-3657</position>
<input>
<ID>J</ID>2655 </input>
<output>
<ID>Q</ID>2177 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2370</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-909,-3703.5</position>
<input>
<ID>J</ID>2641 </input>
<output>
<ID>Q</ID>2642 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2651 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2371</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-916,-3695</position>
<input>
<ID>J</ID>2643 </input>
<output>
<ID>Q</ID>2644 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2651 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2372</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-925,-3687</position>
<input>
<ID>J</ID>2645 </input>
<output>
<ID>Q</ID>2646 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2651 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2373</ID>
<type>AA_AND2</type>
<position>-781,-3661.5</position>
<input>
<ID>IN_0</ID>2177 </input>
<input>
<ID>IN_1</ID>2544 </input>
<output>
<ID>OUT</ID>2679 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2374</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-932,-3678.5</position>
<input>
<ID>J</ID>2647 </input>
<output>
<ID>Q</ID>2648 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2651 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2375</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-940,-3670</position>
<input>
<ID>J</ID>2649 </input>
<output>
<ID>Q</ID>2650 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2651 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2376</ID>
<type>AA_AND2</type>
<position>-782,-3712</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2679 </input>
<output>
<ID>OUT</ID>2680 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2377</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-869.5,-4445.5</position>
<input>
<ID>J</ID>2546 </input>
<output>
<ID>Q</ID>2547 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2571 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2378</ID>
<type>AA_AND2</type>
<position>-768.5,-3709</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2679 </input>
<output>
<ID>OUT</ID>2681 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2379</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-882.5,-4435.5</position>
<input>
<ID>J</ID>2548 </input>
<output>
<ID>Q</ID>2549 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2571 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2380</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-895.5,-4424.5</position>
<input>
<ID>J</ID>2550 </input>
<output>
<ID>Q</ID>2551 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2571 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2381</ID>
<type>AA_AND2</type>
<position>-769,-3701.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2679 </input>
<output>
<ID>OUT</ID>2682 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2382</ID>
<type>AI_XOR2</type>
<position>-792,-4530.5</position>
<input>
<ID>IN_0</ID>2543 </input>
<input>
<ID>IN_1</ID>2545 </input>
<output>
<ID>OUT</ID>2166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2383</ID>
<type>AA_AND2</type>
<position>-768,-3693.5</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2679 </input>
<output>
<ID>OUT</ID>2683 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2384</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-903,-4415.5</position>
<input>
<ID>J</ID>2565 </input>
<output>
<ID>Q</ID>2566 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2571 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2385</ID>
<type>AA_AND2</type>
<position>-768,-3687.5</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2679 </input>
<output>
<ID>OUT</ID>2684 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2386</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-911.5,-4408</position>
<input>
<ID>J</ID>2567 </input>
<output>
<ID>Q</ID>2568 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2571 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2387</ID>
<type>CC_PULSE</type>
<position>-948,-3658</position>
<output>
<ID>OUT_0</ID>2651 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2388</ID>
<type>AA_AND2</type>
<position>-767.5,-3682</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2679 </input>
<output>
<ID>OUT</ID>2685 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2389</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-920.5,-4400.5</position>
<input>
<ID>J</ID>2569 </input>
<output>
<ID>Q</ID>2570 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2571 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2390</ID>
<type>AI_XOR2</type>
<position>-760,-3765.5</position>
<input>
<ID>IN_0</ID>2686 </input>
<input>
<ID>IN_1</ID>2687 </input>
<output>
<ID>OUT</ID>2688 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2391</ID>
<type>CC_PULSE</type>
<position>-950.5,-3502.5</position>
<output>
<ID>OUT_0</ID>2652 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2392</ID>
<type>CC_PULSE</type>
<position>-928.5,-4392.5</position>
<output>
<ID>OUT_0</ID>2571 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2393</ID>
<type>BA_NAND2</type>
<position>-645.5,-3632.5</position>
<input>
<ID>IN_0</ID>2688 </input>
<input>
<ID>IN_1</ID>2687 </input>
<output>
<ID>OUT</ID>2163 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2394</ID>
<type>AA_AND2</type>
<position>-934.5,-4443.5</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2395</ID>
<type>AA_TOGGLE</type>
<position>-787.5,-3478.5</position>
<output>
<ID>OUT_0</ID>2653 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2396</ID>
<type>AA_AND2</type>
<position>-935,-4433.5</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2548 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2397</ID>
<type>AA_AND2</type>
<position>-936.5,-4422.5</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2550 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2398</ID>
<type>AA_AND2</type>
<position>-937,-4413.5</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2565 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2399</ID>
<type>AA_AND2</type>
<position>-938,-4406</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2567 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2400</ID>
<type>AA_AND2</type>
<position>-939,-4398.5</position>
<input>
<ID>IN_0</ID>2387 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2569 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2401</ID>
<type>AE_DFF_LOW</type>
<position>-844.5,-4491</position>
<input>
<ID>IN_0</ID>2388 </input>
<output>
<ID>OUT_0</ID>2395 </output>
<input>
<ID>clear</ID>2256 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2402</ID>
<type>AE_DFF_LOW</type>
<position>-826.5,-4725.5</position>
<input>
<ID>IN_0</ID>2574 </input>
<output>
<ID>OUT_0</ID>2580 </output>
<input>
<ID>clear</ID>2261 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2403</ID>
<type>AE_DFF_LOW</type>
<position>-813,-4725.5</position>
<input>
<ID>IN_0</ID>2575 </input>
<output>
<ID>OUT_0</ID>2581 </output>
<input>
<ID>clear</ID>2261 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2404</ID>
<type>AE_DFF_LOW</type>
<position>-798,-4725.5</position>
<input>
<ID>IN_0</ID>2576 </input>
<output>
<ID>OUT_0</ID>2582 </output>
<input>
<ID>clear</ID>2261 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2405</ID>
<type>AE_DFF_LOW</type>
<position>-787.5,-4725.5</position>
<input>
<ID>IN_0</ID>2577 </input>
<output>
<ID>OUT_0</ID>2583 </output>
<input>
<ID>clear</ID>2261 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2406</ID>
<type>AE_DFF_LOW</type>
<position>-774.5,-4725.5</position>
<input>
<ID>IN_0</ID>2578 </input>
<output>
<ID>OUT_0</ID>2584 </output>
<input>
<ID>clear</ID>2261 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2407</ID>
<type>AE_SMALL_INVERTER</type>
<position>-835.5,-4733</position>
<input>
<ID>IN_0</ID>2579 </input>
<output>
<ID>OUT_0</ID>2585 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2408</ID>
<type>AE_SMALL_INVERTER</type>
<position>-820.5,-4733</position>
<input>
<ID>IN_0</ID>2580 </input>
<output>
<ID>OUT_0</ID>2586 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2409</ID>
<type>AE_SMALL_INVERTER</type>
<position>-805.5,-4733</position>
<input>
<ID>IN_0</ID>2581 </input>
<output>
<ID>OUT_0</ID>2587 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2410</ID>
<type>AE_SMALL_INVERTER</type>
<position>-794,-4732.5</position>
<input>
<ID>IN_0</ID>2582 </input>
<output>
<ID>OUT_0</ID>2588 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2411</ID>
<type>AE_SMALL_INVERTER</type>
<position>-781,-4733</position>
<input>
<ID>IN_0</ID>2583 </input>
<output>
<ID>OUT_0</ID>2589 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2412</ID>
<type>AE_SMALL_INVERTER</type>
<position>-768,-4732.5</position>
<input>
<ID>IN_0</ID>2584 </input>
<output>
<ID>OUT_0</ID>2590 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2413</ID>
<type>AA_AND4</type>
<position>-817.5,-4749.5</position>
<input>
<ID>IN_0</ID>2588 </input>
<input>
<ID>IN_1</ID>2587 </input>
<input>
<ID>IN_2</ID>2586 </input>
<input>
<ID>IN_3</ID>2585 </input>
<output>
<ID>OUT</ID>2591 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2414</ID>
<type>AA_LABEL</type>
<position>-927,-4619</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2415</ID>
<type>AA_AND2</type>
<position>-781,-4748.5</position>
<input>
<ID>IN_0</ID>2590 </input>
<input>
<ID>IN_1</ID>2589 </input>
<output>
<ID>OUT</ID>2592 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2416</ID>
<type>AA_AND2</type>
<position>-803.5,-4771.5</position>
<input>
<ID>IN_0</ID>2592 </input>
<input>
<ID>IN_1</ID>2591 </input>
<output>
<ID>OUT</ID>2316 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2417</ID>
<type>AI_XOR2</type>
<position>-846.5,-4716.5</position>
<input>
<ID>IN_0</ID>2309 </input>
<input>
<ID>IN_1</ID>2594 </input>
<output>
<ID>OUT</ID>2573 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2418</ID>
<type>AI_XOR2</type>
<position>-833,-4716.5</position>
<input>
<ID>IN_0</ID>2311 </input>
<input>
<ID>IN_1</ID>2596 </input>
<output>
<ID>OUT</ID>2574 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2419</ID>
<type>AI_XOR2</type>
<position>-820,-4716.5</position>
<input>
<ID>IN_0</ID>2660 </input>
<input>
<ID>IN_1</ID>2598 </input>
<output>
<ID>OUT</ID>2575 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2420</ID>
<type>AI_XOR2</type>
<position>-807,-4716.5</position>
<input>
<ID>IN_0</ID>2312 </input>
<input>
<ID>IN_1</ID>2600 </input>
<output>
<ID>OUT</ID>2576 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2421</ID>
<type>AI_XOR2</type>
<position>-794.5,-4717</position>
<input>
<ID>IN_0</ID>2313 </input>
<input>
<ID>IN_1</ID>2602 </input>
<output>
<ID>OUT</ID>2577 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2422</ID>
<type>BA_NAND2</type>
<position>-555.5,-3634</position>
<input>
<ID>IN_0</ID>2329 </input>
<input>
<ID>IN_1</ID>2328 </input>
<output>
<ID>OUT</ID>2333 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2423</ID>
<type>AI_XOR2</type>
<position>-782,-4717</position>
<input>
<ID>IN_0</ID>2314 </input>
<input>
<ID>IN_1</ID>2604 </input>
<output>
<ID>OUT</ID>2578 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2424</ID>
<type>AA_LABEL</type>
<position>-980,-4595</position>
<gparam>LABEL_TEXT Zone 7</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2425</ID>
<type>AA_AND4</type>
<position>-575.5,-3615</position>
<input>
<ID>IN_0</ID>2330 </input>
<input>
<ID>IN_1</ID>2331 </input>
<input>
<ID>IN_2</ID>2332 </input>
<input>
<ID>IN_3</ID>2333 </input>
<output>
<ID>OUT</ID>2335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2426</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-867.5,-4679.5</position>
<input>
<ID>J</ID>2593 </input>
<output>
<ID>Q</ID>2594 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2605 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2427</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-880.5,-4669.5</position>
<input>
<ID>J</ID>2595 </input>
<output>
<ID>Q</ID>2596 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2605 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2428</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-893.5,-4658.5</position>
<input>
<ID>J</ID>2597 </input>
<output>
<ID>Q</ID>2598 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2605 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2429</ID>
<type>AI_XOR2</type>
<position>-790,-4764.5</position>
<input>
<ID>IN_0</ID>2591 </input>
<input>
<ID>IN_1</ID>2592 </input>
<output>
<ID>OUT</ID>2168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2430</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-901,-4649.5</position>
<input>
<ID>J</ID>2599 </input>
<output>
<ID>Q</ID>2600 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2605 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2431</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-909.5,-4642</position>
<input>
<ID>J</ID>2601 </input>
<output>
<ID>Q</ID>2602 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2605 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2432</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-918.5,-4634.5</position>
<input>
<ID>J</ID>2603 </input>
<output>
<ID>Q</ID>2604 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2605 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2433</ID>
<type>CC_PULSE</type>
<position>-926.5,-4626.5</position>
<output>
<ID>OUT_0</ID>2605 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2434</ID>
<type>AA_AND2</type>
<position>-932.5,-4677.5</position>
<input>
<ID>IN_0</ID>2572 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2435</ID>
<type>AA_AND2</type>
<position>-933,-4667.5</position>
<input>
<ID>IN_0</ID>2572 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2436</ID>
<type>AA_AND2</type>
<position>-934.5,-4656.5</position>
<input>
<ID>IN_0</ID>2572 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2437</ID>
<type>AA_AND2</type>
<position>-935,-4647.5</position>
<input>
<ID>IN_0</ID>2572 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2438</ID>
<type>AA_AND2</type>
<position>-936,-4640</position>
<input>
<ID>IN_0</ID>2572 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2439</ID>
<type>AA_AND2</type>
<position>-937,-4632.5</position>
<input>
<ID>IN_0</ID>2572 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2603 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2440</ID>
<type>AE_DFF_LOW</type>
<position>-842.5,-4725</position>
<input>
<ID>IN_0</ID>2573 </input>
<output>
<ID>OUT_0</ID>2579 </output>
<input>
<ID>clear</ID>2261 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2441</ID>
<type>AE_DFF_LOW</type>
<position>-817.5,-4952.5</position>
<input>
<ID>IN_0</ID>2608 </input>
<output>
<ID>OUT_0</ID>2614 </output>
<input>
<ID>clear</ID>2659 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2442</ID>
<type>AE_DFF_LOW</type>
<position>-804,-4952.5</position>
<input>
<ID>IN_0</ID>2609 </input>
<output>
<ID>OUT_0</ID>2615 </output>
<input>
<ID>clear</ID>2659 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2443</ID>
<type>AE_DFF_LOW</type>
<position>-789,-4952.5</position>
<input>
<ID>IN_0</ID>2610 </input>
<output>
<ID>OUT_0</ID>2616 </output>
<input>
<ID>clear</ID>2659 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2444</ID>
<type>AE_DFF_LOW</type>
<position>-778.5,-4952.5</position>
<input>
<ID>IN_0</ID>2611 </input>
<output>
<ID>OUT_0</ID>2617 </output>
<input>
<ID>clear</ID>2659 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2445</ID>
<type>AE_DFF_LOW</type>
<position>-765.5,-4952.5</position>
<input>
<ID>IN_0</ID>2612 </input>
<output>
<ID>OUT_0</ID>2618 </output>
<input>
<ID>clear</ID>2659 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2446</ID>
<type>AE_SMALL_INVERTER</type>
<position>-826.5,-4960</position>
<input>
<ID>IN_0</ID>2613 </input>
<output>
<ID>OUT_0</ID>2619 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2447</ID>
<type>AE_SMALL_INVERTER</type>
<position>-811.5,-4960</position>
<input>
<ID>IN_0</ID>2614 </input>
<output>
<ID>OUT_0</ID>2620 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2448</ID>
<type>AE_SMALL_INVERTER</type>
<position>-796.5,-4960</position>
<input>
<ID>IN_0</ID>2615 </input>
<output>
<ID>OUT_0</ID>2621 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2449</ID>
<type>AE_SMALL_INVERTER</type>
<position>-785,-4959.5</position>
<input>
<ID>IN_0</ID>2616 </input>
<output>
<ID>OUT_0</ID>2622 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2450</ID>
<type>AE_SMALL_INVERTER</type>
<position>-772,-4960</position>
<input>
<ID>IN_0</ID>2617 </input>
<output>
<ID>OUT_0</ID>2623 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2451</ID>
<type>AE_SMALL_INVERTER</type>
<position>-759,-4959.5</position>
<input>
<ID>IN_0</ID>2618 </input>
<output>
<ID>OUT_0</ID>2624 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2452</ID>
<type>AA_AND4</type>
<position>-808.5,-4976.5</position>
<input>
<ID>IN_0</ID>2622 </input>
<input>
<ID>IN_1</ID>2621 </input>
<input>
<ID>IN_2</ID>2620 </input>
<input>
<ID>IN_3</ID>2619 </input>
<output>
<ID>OUT</ID>2625 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2453</ID>
<type>AA_LABEL</type>
<position>-918,-4846</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2454</ID>
<type>AA_AND2</type>
<position>-772,-4975.5</position>
<input>
<ID>IN_0</ID>2624 </input>
<input>
<ID>IN_1</ID>2623 </input>
<output>
<ID>OUT</ID>2626 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2455</ID>
<type>AA_AND2</type>
<position>-794.5,-4998.5</position>
<input>
<ID>IN_0</ID>2626 </input>
<input>
<ID>IN_1</ID>2625 </input>
<output>
<ID>OUT</ID>2328 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2456</ID>
<type>AI_XOR2</type>
<position>-837.5,-4943.5</position>
<input>
<ID>IN_0</ID>2319 </input>
<input>
<ID>IN_1</ID>2628 </input>
<output>
<ID>OUT</ID>2607 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2457</ID>
<type>AI_XOR2</type>
<position>-824,-4943.5</position>
<input>
<ID>IN_0</ID>2321 </input>
<input>
<ID>IN_1</ID>2630 </input>
<output>
<ID>OUT</ID>2608 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2458</ID>
<type>AI_XOR2</type>
<position>-811,-4943.5</position>
<input>
<ID>IN_0</ID>2322 </input>
<input>
<ID>IN_1</ID>2632 </input>
<output>
<ID>OUT</ID>2609 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2459</ID>
<type>AI_XOR2</type>
<position>-798,-4943.5</position>
<input>
<ID>IN_0</ID>2323 </input>
<input>
<ID>IN_1</ID>2634 </input>
<output>
<ID>OUT</ID>2610 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2460</ID>
<type>AI_XOR2</type>
<position>-785.5,-4944</position>
<input>
<ID>IN_0</ID>2324 </input>
<input>
<ID>IN_1</ID>2636 </input>
<output>
<ID>OUT</ID>2611 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2461</ID>
<type>AI_XOR2</type>
<position>-773,-4944</position>
<input>
<ID>IN_0</ID>2325 </input>
<input>
<ID>IN_1</ID>2638 </input>
<output>
<ID>OUT</ID>2612 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2462</ID>
<type>AA_AND2</type>
<position>-613.5,-3593</position>
<input>
<ID>IN_0</ID>2334 </input>
<input>
<ID>IN_1</ID>2335 </input>
<output>
<ID>OUT</ID>2348 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2463</ID>
<type>AA_LABEL</type>
<position>-975,-4809</position>
<gparam>LABEL_TEXT Zone 8</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2464</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-858.5,-4906.5</position>
<input>
<ID>J</ID>2627 </input>
<output>
<ID>Q</ID>2628 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2639 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2465</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-871.5,-4896.5</position>
<input>
<ID>J</ID>2629 </input>
<output>
<ID>Q</ID>2630 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2639 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2466</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-884.5,-4885.5</position>
<input>
<ID>J</ID>2631 </input>
<output>
<ID>Q</ID>2632 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2639 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2467</ID>
<type>AI_XOR2</type>
<position>-781,-4991.5</position>
<input>
<ID>IN_0</ID>2625 </input>
<input>
<ID>IN_1</ID>2626 </input>
<output>
<ID>OUT</ID>2170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2468</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-892,-4876.5</position>
<input>
<ID>J</ID>2633 </input>
<output>
<ID>Q</ID>2634 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2639 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2469</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-900.5,-4869</position>
<input>
<ID>J</ID>2635 </input>
<output>
<ID>Q</ID>2636 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2639 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2470</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-909.5,-4861.5</position>
<input>
<ID>J</ID>2637 </input>
<output>
<ID>Q</ID>2638 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2639 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2471</ID>
<type>CC_PULSE</type>
<position>-917.5,-4853.5</position>
<output>
<ID>OUT_0</ID>2639 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2472</ID>
<type>AA_AND2</type>
<position>-923.5,-4904.5</position>
<input>
<ID>IN_0</ID>2606 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2473</ID>
<type>AA_AND2</type>
<position>-924,-4894.5</position>
<input>
<ID>IN_0</ID>2606 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2629 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2474</ID>
<type>AA_AND2</type>
<position>-925.5,-4883.5</position>
<input>
<ID>IN_0</ID>2606 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2631 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2475</ID>
<type>AA_AND2</type>
<position>-926,-4874.5</position>
<input>
<ID>IN_0</ID>2606 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2633 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2476</ID>
<type>AA_AND2</type>
<position>-927,-4867</position>
<input>
<ID>IN_0</ID>2606 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2635 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2477</ID>
<type>AA_AND2</type>
<position>-928,-4859.5</position>
<input>
<ID>IN_0</ID>2606 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2637 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2478</ID>
<type>AE_DFF_LOW</type>
<position>-833.5,-4952</position>
<input>
<ID>IN_0</ID>2607 </input>
<output>
<ID>OUT_0</ID>2613 </output>
<input>
<ID>clear</ID>2659 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2479</ID>
<type>AA_LABEL</type>
<position>-795,-3471.5</position>
<gparam>LABEL_TEXT Reset Storage before saving</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2480</ID>
<type>AA_LABEL</type>
<position>-873.5,-3785</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2482</ID>
<type>AA_LABEL</type>
<position>-1312,-3181.5</position>
<gparam>LABEL_TEXT Insert values first to start the counter</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2484</ID>
<type>AA_LABEL</type>
<position>-883,-3326</position>
<gparam>LABEL_TEXT Minutes Output</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2486</ID>
<type>AA_LABEL</type>
<position>-1299.5,-3610</position>
<gparam>LABEL_TEXT Timer Output</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2488</ID>
<type>AA_LABEL</type>
<position>-781,-3593.5</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2489</ID>
<type>AA_LABEL</type>
<position>-778.5,-3716</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2490</ID>
<type>AA_LABEL</type>
<position>-774,-3876</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2491</ID>
<type>AA_LABEL</type>
<position>-764,-4062.5</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2492</ID>
<type>AA_LABEL</type>
<position>-753,-4261</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2493</ID>
<type>AA_LABEL</type>
<position>-760.5,-4480</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2494</ID>
<type>AA_LABEL</type>
<position>-748,-4715</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2495</ID>
<type>AA_LABEL</type>
<position>-739,-4943</position>
<gparam>LABEL_TEXT Values being compared</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2497</ID>
<type>AA_LABEL</type>
<position>-500.5,-3607.5</position>
<gparam>LABEL_TEXT Conditions to reset timer when particular zone finishes watering</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2499</ID>
<type>AA_LABEL</type>
<position>-763.5,-3568</position>
<gparam>LABEL_TEXT Minutes Output</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2500</ID>
<type>AA_LABEL</type>
<position>-676.5,-3692.5</position>
<gparam>LABEL_TEXT Minutes Output</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2502</ID>
<type>AA_LABEL</type>
<position>-731.5,-3670</position>
<gparam>LABEL_TEXT Conditions being checked it that particular zone is selected and the previous zone is finished.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1860</ID>
<type>AE_DFF_LOW</type>
<position>-840.5,-3888.5</position>
<input>
<ID>IN_0</ID>2205 </input>
<output>
<ID>OUT_0</ID>2213 </output>
<input>
<ID>clear</ID>2678 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1861</ID>
<type>AE_OR2</type>
<position>-790.5,-3647</position>
<input>
<ID>IN_0</ID>2156 </input>
<input>
<ID>IN_1</ID>2393 </input>
<output>
<ID>OUT</ID>2654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1862</ID>
<type>AA_LABEL</type>
<position>-920,-3470</position>
<gparam>LABEL_TEXT Keep Off before setting value and then turn it on</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1863</ID>
<type>AE_OR2</type>
<position>-789.5,-3931</position>
<input>
<ID>IN_0</ID>2158 </input>
<input>
<ID>IN_1</ID>2174 </input>
<output>
<ID>OUT</ID>2183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1864</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-808.5,-3774</position>
<input>
<ID>J</ID>2687 </input>
<output>
<ID>Q</ID>2157 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1865</ID>
<type>AI_XOR2</type>
<position>-785.5,-3757.5</position>
<input>
<ID>IN_0</ID>2386 </input>
<input>
<ID>IN_1</ID>2385 </input>
<output>
<ID>OUT</ID>2160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1866</ID>
<type>AA_AND4</type>
<position>-640.5,-3616.5</position>
<input>
<ID>IN_0</ID>2159 </input>
<input>
<ID>IN_1</ID>2163 </input>
<input>
<ID>IN_2</ID>2180 </input>
<input>
<ID>IN_3</ID>2181 </input>
<output>
<ID>OUT</ID>2334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1867</ID>
<type>AE_OR2</type>
<position>-771.5,-3764</position>
<input>
<ID>IN_0</ID>2160 </input>
<input>
<ID>IN_1</ID>2544 </input>
<output>
<ID>OUT</ID>2686 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1868</ID>
<type>AA_AND2</type>
<position>-788.5,-3779</position>
<input>
<ID>IN_0</ID>2157 </input>
<input>
<ID>IN_1</ID>2174 </input>
<output>
<ID>OUT</ID>2161 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1869</ID>
<type>GA_LED</type>
<position>-747.5,-3764</position>
<input>
<ID>N_in0</ID>2688 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1870</ID>
<type>AE_DFF_LOW</type>
<position>-827,-3888.5</position>
<input>
<ID>IN_0</ID>2206 </input>
<output>
<ID>OUT_0</ID>2214 </output>
<input>
<ID>clear</ID>2678 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1871</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-919.5,-4081.5</position>
<input>
<ID>J</ID>2167 </input>
<output>
<ID>Q</ID>2246 </output>
<input>
<ID>clear</ID>2167 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2169 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1872</ID>
<type>AA_AND2</type>
<position>-930,-4091.5</position>
<input>
<ID>IN_0</ID>2303 </input>
<input>
<ID>IN_1</ID>2182 </input>
<output>
<ID>OUT</ID>2165 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1873</ID>
<type>AA_AND2</type>
<position>-780.5,-3861</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2161 </input>
<output>
<ID>OUT</ID>2171 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1874</ID>
<type>AE_OR2</type>
<position>-783,-4110.5</position>
<input>
<ID>IN_0</ID>2162 </input>
<input>
<ID>IN_1</ID>2279 </input>
<output>
<ID>OUT</ID>2230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1875</ID>
<type>AE_SMALL_INVERTER</type>
<position>-937.5,-4087.5</position>
<input>
<ID>IN_0</ID>2165 </input>
<output>
<ID>OUT_0</ID>2167 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1876</ID>
<type>AE_OR2</type>
<position>-775,-4309.5</position>
<input>
<ID>IN_0</ID>2164 </input>
<input>
<ID>IN_1</ID>2349 </input>
<output>
<ID>OUT</ID>2273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1877</ID>
<type>AA_AND2</type>
<position>-765,-3855.5</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2161 </input>
<output>
<ID>OUT</ID>2172 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1878</ID>
<type>GA_LED</type>
<position>-752.5,-4531.5</position>
<input>
<ID>N_in0</ID>2307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1879</ID>
<type>GA_LED</type>
<position>-912.5,-4083.5</position>
<input>
<ID>N_in0</ID>2169 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1880</ID>
<type>AE_OR2</type>
<position>-779.5,-4531.5</position>
<input>
<ID>IN_0</ID>2166 </input>
<input>
<ID>IN_1</ID>2387 </input>
<output>
<ID>OUT</ID>2305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1881</ID>
<type>AE_DFF_LOW</type>
<position>-812,-3888.5</position>
<input>
<ID>IN_0</ID>2209 </input>
<output>
<ID>OUT_0</ID>2215 </output>
<input>
<ID>clear</ID>2678 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1882</ID>
<type>AA_AND2</type>
<position>-764.5,-3847.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2161 </input>
<output>
<ID>OUT</ID>2173 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1883</ID>
<type>AE_OR2</type>
<position>-778,-4765.5</position>
<input>
<ID>IN_0</ID>2168 </input>
<input>
<ID>IN_1</ID>2572 </input>
<output>
<ID>OUT</ID>2315 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1884</ID>
<type>AE_DFF_LOW</type>
<position>-801.5,-3888.5</position>
<input>
<ID>IN_0</ID>2210 </input>
<output>
<ID>OUT_0</ID>2216 </output>
<input>
<ID>clear</ID>2678 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1885</ID>
<type>AE_DFF_LOW</type>
<position>-788.5,-3888.5</position>
<input>
<ID>IN_0</ID>2211 </input>
<output>
<ID>OUT_0</ID>2217 </output>
<input>
<ID>clear</ID>2678 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1886</ID>
<type>GA_LED</type>
<position>-755,-4765</position>
<input>
<ID>N_in0</ID>2317 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1887</ID>
<type>AA_AND2</type>
<position>-763.5,-3839.5</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2161 </input>
<output>
<ID>OUT</ID>2175 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1888</ID>
<type>AA_AND2</type>
<position>-889.5,-4089.5</position>
<input>
<ID>IN_0</ID>2298 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2182 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1889</ID>
<type>AA_AND2</type>
<position>-763,-3829</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2161 </input>
<output>
<ID>OUT</ID>2176 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1890</ID>
<type>AE_SMALL_INVERTER</type>
<position>-849.5,-3896</position>
<input>
<ID>IN_0</ID>2212 </input>
<output>
<ID>OUT_0</ID>2218 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1891</ID>
<type>GA_LED</type>
<position>-740,-4993</position>
<input>
<ID>N_in0</ID>2329 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1892</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-901.5,-4290</position>
<input>
<ID>J</ID>2248 </input>
<output>
<ID>Q</ID>2251 </output>
<input>
<ID>clear</ID>2248 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2249 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1893</ID>
<type>AE_OR2</type>
<position>-769,-4992.5</position>
<input>
<ID>IN_0</ID>2170 </input>
<input>
<ID>IN_1</ID>2606 </input>
<output>
<ID>OUT</ID>2326 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1894</ID>
<type>AA_AND2</type>
<position>-763.5,-3818</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2161 </input>
<output>
<ID>OUT</ID>2178 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1895</ID>
<type>AA_AND2</type>
<position>-912,-4300</position>
<input>
<ID>IN_0</ID>2369 </input>
<input>
<ID>IN_1</ID>2250 </input>
<output>
<ID>OUT</ID>2247 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1896</ID>
<type>BA_NAND2</type>
<position>-626,-3632.5</position>
<input>
<ID>IN_0</ID>2184 </input>
<input>
<ID>IN_1</ID>2179 </input>
<output>
<ID>OUT</ID>2180 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1897</ID>
<type>AE_SMALL_INVERTER</type>
<position>-919.5,-4296</position>
<input>
<ID>IN_0</ID>2247 </input>
<output>
<ID>OUT_0</ID>2248 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1898</ID>
<type>GA_LED</type>
<position>-894.5,-4292</position>
<input>
<ID>N_in0</ID>2249 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1899</ID>
<type>AE_SMALL_INVERTER</type>
<position>-834.5,-3896</position>
<input>
<ID>IN_0</ID>2213 </input>
<output>
<ID>OUT_0</ID>2219 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1900</ID>
<type>AI_XOR2</type>
<position>-776.5,-3932</position>
<input>
<ID>IN_0</ID>2183 </input>
<input>
<ID>IN_1</ID>2179 </input>
<output>
<ID>OUT</ID>2184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1901</ID>
<type>AA_AND2</type>
<position>-871.5,-4298</position>
<input>
<ID>IN_0</ID>2368 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2250 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1902</ID>
<type>GA_LED</type>
<position>-758.5,-3926</position>
<input>
<ID>N_in0</ID>2184 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1903</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-903,-4513</position>
<input>
<ID>J</ID>2253 </input>
<output>
<ID>Q</ID>2256 </output>
<input>
<ID>clear</ID>2253 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2254 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1904</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-802.5,-3943</position>
<input>
<ID>J</ID>2179 </input>
<output>
<ID>Q</ID>2201 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1905</ID>
<type>AE_SMALL_INVERTER</type>
<position>-819.5,-3896</position>
<input>
<ID>IN_0</ID>2214 </input>
<output>
<ID>OUT_0</ID>2221 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1906</ID>
<type>AA_AND2</type>
<position>-913.5,-4523</position>
<input>
<ID>IN_0</ID>2545 </input>
<input>
<ID>IN_1</ID>2255 </input>
<output>
<ID>OUT</ID>2252 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1907</ID>
<type>AE_SMALL_INVERTER</type>
<position>-808,-3895.5</position>
<input>
<ID>IN_0</ID>2215 </input>
<output>
<ID>OUT_0</ID>2222 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1908</ID>
<type>AA_TOGGLE</type>
<position>-994.5,-3490.5</position>
<output>
<ID>OUT_0</ID>2689 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1909</ID>
<type>AA_LABEL</type>
<position>-946,-3652.5</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1910</ID>
<type>AA_LABEL</type>
<position>-950.5,-3495</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1911</ID>
<type>AE_SMALL_INVERTER</type>
<position>-795,-3896</position>
<input>
<ID>IN_0</ID>2216 </input>
<output>
<ID>OUT_0</ID>2224 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1912</ID>
<type>AE_SMALL_INVERTER</type>
<position>-782,-3895.5</position>
<input>
<ID>IN_0</ID>2217 </input>
<output>
<ID>OUT_0</ID>2225 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1913</ID>
<type>AI_XOR2</type>
<position>-775.5,-3647.5</position>
<input>
<ID>IN_0</ID>2654 </input>
<input>
<ID>IN_1</ID>2655 </input>
<output>
<ID>OUT</ID>2656 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1914</ID>
<type>AA_AND4</type>
<position>-831.5,-3912.5</position>
<input>
<ID>IN_0</ID>2222 </input>
<input>
<ID>IN_1</ID>2221 </input>
<input>
<ID>IN_2</ID>2219 </input>
<input>
<ID>IN_3</ID>2218 </input>
<output>
<ID>OUT</ID>2226 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1915</ID>
<type>AE_DFF_LOW</type>
<position>-850.5,-3726.5</position>
<input>
<ID>IN_0</ID>2186 </input>
<output>
<ID>OUT_0</ID>2192 </output>
<input>
<ID>clear</ID>2673 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1916</ID>
<type>BA_NAND2</type>
<position>-659.5,-3632.5</position>
<input>
<ID>IN_0</ID>2656 </input>
<input>
<ID>IN_1</ID>2655 </input>
<output>
<ID>OUT</ID>2159 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1917</ID>
<type>AE_DFF_LOW</type>
<position>-837,-3726.5</position>
<input>
<ID>IN_0</ID>2187 </input>
<output>
<ID>OUT_0</ID>2193 </output>
<input>
<ID>clear</ID>2673 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1918</ID>
<type>AA_LABEL</type>
<position>-941,-3782</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1919</ID>
<type>AE_DFF_LOW</type>
<position>-822,-3726.5</position>
<input>
<ID>IN_0</ID>2188 </input>
<output>
<ID>OUT_0</ID>2194 </output>
<input>
<ID>clear</ID>2673 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1920</ID>
<type>AE_DFF_LOW</type>
<position>-811.5,-3726.5</position>
<input>
<ID>IN_0</ID>2189 </input>
<output>
<ID>OUT_0</ID>2195 </output>
<input>
<ID>clear</ID>2673 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1921</ID>
<type>AE_DFF_LOW</type>
<position>-798.5,-3726.5</position>
<input>
<ID>IN_0</ID>2190 </input>
<output>
<ID>OUT_0</ID>2196 </output>
<input>
<ID>clear</ID>2673 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1922</ID>
<type>AA_AND2</type>
<position>-795,-3911.5</position>
<input>
<ID>IN_0</ID>2225 </input>
<input>
<ID>IN_1</ID>2224 </input>
<output>
<ID>OUT</ID>2227 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1923</ID>
<type>AE_SMALL_INVERTER</type>
<position>-859.5,-3734</position>
<input>
<ID>IN_0</ID>2191 </input>
<output>
<ID>OUT_0</ID>2197 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1924</ID>
<type>AA_AND2</type>
<position>-817.5,-3934.5</position>
<input>
<ID>IN_0</ID>2227 </input>
<input>
<ID>IN_1</ID>2226 </input>
<output>
<ID>OUT</ID>2179 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1925</ID>
<type>AE_SMALL_INVERTER</type>
<position>-844.5,-3734</position>
<input>
<ID>IN_0</ID>2192 </input>
<output>
<ID>OUT_0</ID>2198 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1926</ID>
<type>AE_SMALL_INVERTER</type>
<position>-829.5,-3734</position>
<input>
<ID>IN_0</ID>2193 </input>
<output>
<ID>OUT_0</ID>2199 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1927</ID>
<type>AE_SMALL_INVERTER</type>
<position>-818,-3733.5</position>
<input>
<ID>IN_0</ID>2194 </input>
<output>
<ID>OUT_0</ID>2200 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1928</ID>
<type>AE_SMALL_INVERTER</type>
<position>-805,-3734</position>
<input>
<ID>IN_0</ID>2195 </input>
<output>
<ID>OUT_0</ID>2383 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1929</ID>
<type>AE_SMALL_INVERTER</type>
<position>-792,-3733.5</position>
<input>
<ID>IN_0</ID>2196 </input>
<output>
<ID>OUT_0</ID>2384 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1930</ID>
<type>AI_XOR2</type>
<position>-860.5,-3879.5</position>
<input>
<ID>IN_0</ID>2171 </input>
<input>
<ID>IN_1</ID>2232 </input>
<output>
<ID>OUT</ID>2202 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1931</ID>
<type>AI_XOR2</type>
<position>-847,-3879.5</position>
<input>
<ID>IN_0</ID>2172 </input>
<input>
<ID>IN_1</ID>2234 </input>
<output>
<ID>OUT</ID>2205 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1932</ID>
<type>AI_XOR2</type>
<position>-834,-3879.5</position>
<input>
<ID>IN_0</ID>2173 </input>
<input>
<ID>IN_1</ID>2236 </input>
<output>
<ID>OUT</ID>2206 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1933</ID>
<type>AI_XOR2</type>
<position>-821,-3879.5</position>
<input>
<ID>IN_0</ID>2175 </input>
<input>
<ID>IN_1</ID>2238 </input>
<output>
<ID>OUT</ID>2209 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1934</ID>
<type>AI_XOR2</type>
<position>-808.5,-3880</position>
<input>
<ID>IN_0</ID>2176 </input>
<input>
<ID>IN_1</ID>2240 </input>
<output>
<ID>OUT</ID>2210 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1935</ID>
<type>AA_AND2</type>
<position>-783,-3947</position>
<input>
<ID>IN_0</ID>2201 </input>
<input>
<ID>IN_1</ID>2279 </input>
<output>
<ID>OUT</ID>2204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1936</ID>
<type>AI_XOR2</type>
<position>-796,-3880</position>
<input>
<ID>IN_0</ID>2178 </input>
<input>
<ID>IN_1</ID>2242 </input>
<output>
<ID>OUT</ID>2211 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1937</ID>
<type>AE_SMALL_INVERTER</type>
<position>-921,-4519</position>
<input>
<ID>IN_0</ID>2252 </input>
<output>
<ID>OUT_0</ID>2253 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1938</ID>
<type>AA_LABEL</type>
<position>-1004,-3760</position>
<gparam>LABEL_TEXT Zone 3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1939</ID>
<type>AA_AND2</type>
<position>-778,-4043</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2204 </input>
<output>
<ID>OUT</ID>2203 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1940</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-881.5,-3842.5</position>
<input>
<ID>J</ID>2231 </input>
<output>
<ID>Q</ID>2232 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2243 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1941</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-894.5,-3832.5</position>
<input>
<ID>J</ID>2233 </input>
<output>
<ID>Q</ID>2234 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2243 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1942</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-907.5,-3821.5</position>
<input>
<ID>J</ID>2235 </input>
<output>
<ID>Q</ID>2236 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2243 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1943</ID>
<type>AI_XOR2</type>
<position>-804,-3927.5</position>
<input>
<ID>IN_0</ID>2226 </input>
<input>
<ID>IN_1</ID>2227 </input>
<output>
<ID>OUT</ID>2158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1944</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-915,-3812.5</position>
<input>
<ID>J</ID>2237 </input>
<output>
<ID>Q</ID>2238 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2243 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1945</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-923.5,-3805</position>
<input>
<ID>J</ID>2239 </input>
<output>
<ID>Q</ID>2240 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2243 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1946</ID>
<type>GA_LED</type>
<position>-762.5,-3647</position>
<input>
<ID>N_in0</ID>2656 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1947</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-932.5,-3797.5</position>
<input>
<ID>J</ID>2241 </input>
<output>
<ID>Q</ID>2242 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2243 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1948</ID>
<type>CC_PULSE</type>
<position>-940.5,-3789.5</position>
<output>
<ID>OUT_0</ID>2243 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>1949</ID>
<type>AA_TOGGLE</type>
<position>-874,-3789.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1950</ID>
<type>AA_AND2</type>
<position>-946.5,-3840.5</position>
<input>
<ID>IN_0</ID>2174 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1951</ID>
<type>AA_AND2</type>
<position>-947,-3830.5</position>
<input>
<ID>IN_0</ID>2174 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1952</ID>
<type>AA_AND2</type>
<position>-948.5,-3819.5</position>
<input>
<ID>IN_0</ID>2174 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1953</ID>
<type>AA_AND2</type>
<position>-949,-3810.5</position>
<input>
<ID>IN_0</ID>2174 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1954</ID>
<type>AA_AND2</type>
<position>-950,-3803</position>
<input>
<ID>IN_0</ID>2174 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1955</ID>
<type>AA_AND2</type>
<position>-951,-3795.5</position>
<input>
<ID>IN_0</ID>2174 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1956</ID>
<type>AE_DFF_LOW</type>
<position>-856.5,-3888</position>
<input>
<ID>IN_0</ID>2202 </input>
<output>
<ID>OUT_0</ID>2212 </output>
<input>
<ID>clear</ID>2678 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1957</ID>
<type>GA_LED</type>
<position>-896,-4515</position>
<input>
<ID>N_in0</ID>2254 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1958</ID>
<type>AA_AND2</type>
<position>-768,-4031</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2204 </input>
<output>
<ID>OUT</ID>2207 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1959</ID>
<type>AA_AND2</type>
<position>-768,-4022.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2204 </input>
<output>
<ID>OUT</ID>2220 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1960</ID>
<type>AA_AND2</type>
<position>-873,-4521</position>
<input>
<ID>IN_0</ID>2543 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2255 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1961</ID>
<type>AI_XOR2</type>
<position>-813.5,-3640.5</position>
<input>
<ID>IN_0</ID>2414 </input>
<input>
<ID>IN_1</ID>2415 </input>
<output>
<ID>OUT</ID>2156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1962</ID>
<type>AA_AND2</type>
<position>-767,-4015</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2204 </input>
<output>
<ID>OUT</ID>2223 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1963</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-901,-4746.5</position>
<input>
<ID>J</ID>2258 </input>
<output>
<ID>Q</ID>2261 </output>
<input>
<ID>clear</ID>2258 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2259 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1964</ID>
<type>AA_AND2</type>
<position>-766.5,-4006</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2204 </input>
<output>
<ID>OUT</ID>2228 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1965</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-794.5,-4128.5</position>
<input>
<ID>J</ID>2244 </input>
<output>
<ID>Q</ID>2265 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1966</ID>
<type>AA_AND2</type>
<position>-766,-3998</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2204 </input>
<output>
<ID>OUT</ID>2229 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1967</ID>
<type>AA_AND2</type>
<position>-911.5,-4756.5</position>
<input>
<ID>IN_0</ID>2592 </input>
<input>
<ID>IN_1</ID>2260 </input>
<output>
<ID>OUT</ID>2257 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1968</ID>
<type>AI_XOR2</type>
<position>-768.5,-4111</position>
<input>
<ID>IN_0</ID>2230 </input>
<input>
<ID>IN_1</ID>2244 </input>
<output>
<ID>OUT</ID>2245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1969</ID>
<type>AA_AND2</type>
<position>-785,-4138</position>
<input>
<ID>IN_0</ID>2265 </input>
<input>
<ID>IN_1</ID>2349 </input>
<output>
<ID>OUT</ID>2267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1970</ID>
<type>GA_LED</type>
<position>-748,-4111</position>
<input>
<ID>N_in0</ID>2245 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1971</ID>
<type>AE_SMALL_INVERTER</type>
<position>-919,-4752.5</position>
<input>
<ID>IN_0</ID>2257 </input>
<output>
<ID>OUT_0</ID>2258 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1972</ID>
<type>BA_NAND2</type>
<position>-609.5,-3633</position>
<input>
<ID>IN_0</ID>2245 </input>
<input>
<ID>IN_1</ID>2244 </input>
<output>
<ID>OUT</ID>2181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1973</ID>
<type>AA_AND2</type>
<position>-765.5,-4209.5</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2267 </input>
<output>
<ID>OUT</ID>2266 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1974</ID>
<type>GA_LED</type>
<position>-894,-4748.5</position>
<input>
<ID>N_in0</ID>2259 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1975</ID>
<type>AA_AND2</type>
<position>-753.5,-4201</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2267 </input>
<output>
<ID>OUT</ID>2268 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1976</ID>
<type>AA_AND2</type>
<position>-753.5,-4191</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2267 </input>
<output>
<ID>OUT</ID>2269 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1977</ID>
<type>AA_AND2</type>
<position>-871,-4754.5</position>
<input>
<ID>IN_0</ID>2591 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2260 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1978</ID>
<type>AA_AND2</type>
<position>-752,-4184</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2267 </input>
<output>
<ID>OUT</ID>2270 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1979</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-878.5,-4975</position>
<input>
<ID>J</ID>2263 </input>
<output>
<ID>Q</ID>2659 </output>
<input>
<ID>clear</ID>2263 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2264 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1980</ID>
<type>AA_AND2</type>
<position>-751.5,-4174.5</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2267 </input>
<output>
<ID>OUT</ID>2271 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1981</ID>
<type>AA_AND2</type>
<position>-889,-4985</position>
<input>
<ID>IN_0</ID>2626 </input>
<input>
<ID>IN_1</ID>2658 </input>
<output>
<ID>OUT</ID>2262 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1982</ID>
<type>AA_AND2</type>
<position>-751,-4167.5</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2267 </input>
<output>
<ID>OUT</ID>2272 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1983</ID>
<type>AE_SMALL_INVERTER</type>
<position>-896.5,-4981</position>
<input>
<ID>IN_0</ID>2262 </input>
<output>
<ID>OUT_0</ID>2263 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1984</ID>
<type>AI_XOR2</type>
<position>-763.5,-4310</position>
<input>
<ID>IN_0</ID>2273 </input>
<input>
<ID>IN_1</ID>2274 </input>
<output>
<ID>OUT</ID>2275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1985</ID>
<type>GA_LED</type>
<position>-871.5,-4977</position>
<input>
<ID>N_in0</ID>2264 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1986</ID>
<type>GA_LED</type>
<position>-749.5,-4309.5</position>
<input>
<ID>N_in0</ID>2275 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1987</ID>
<type>BA_NAND2</type>
<position>-594.5,-3633.5</position>
<input>
<ID>IN_0</ID>2275 </input>
<input>
<ID>IN_1</ID>2274 </input>
<output>
<ID>OUT</ID>2330 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1988</ID>
<type>AA_AND2</type>
<position>-848.5,-4983</position>
<input>
<ID>IN_0</ID>2625 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2658 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1989</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-786.5,-4325</position>
<input>
<ID>J</ID>2274 </input>
<output>
<ID>Q</ID>2276 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1990</ID>
<type>AA_AND2</type>
<position>-772,-4333.5</position>
<input>
<ID>IN_0</ID>2276 </input>
<input>
<ID>IN_1</ID>2387 </input>
<output>
<ID>OUT</ID>2277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1991</ID>
<type>AA_AND2</type>
<position>-774.5,-4468</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2277 </input>
<output>
<ID>OUT</ID>2278 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1992</ID>
<type>AA_AND2</type>
<position>-763.5,-4462</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2277 </input>
<output>
<ID>OUT</ID>2299 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1993</ID>
<type>AE_DFF_LOW</type>
<position>-832.5,-4070.5</position>
<input>
<ID>IN_0</ID>2281 </input>
<output>
<ID>OUT_0</ID>2287 </output>
<input>
<ID>clear</ID>2246 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1994</ID>
<type>AE_DFF_LOW</type>
<position>-819,-4070.5</position>
<input>
<ID>IN_0</ID>2282 </input>
<output>
<ID>OUT_0</ID>2288 </output>
<input>
<ID>clear</ID>2246 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1995</ID>
<type>AE_DFF_LOW</type>
<position>-804,-4070.5</position>
<input>
<ID>IN_0</ID>2283 </input>
<output>
<ID>OUT_0</ID>2289 </output>
<input>
<ID>clear</ID>2246 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1996</ID>
<type>AE_DFF_LOW</type>
<position>-793.5,-4070.5</position>
<input>
<ID>IN_0</ID>2284 </input>
<output>
<ID>OUT_0</ID>2290 </output>
<input>
<ID>clear</ID>2246 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1997</ID>
<type>AE_DFF_LOW</type>
<position>-780.5,-4070.5</position>
<input>
<ID>IN_0</ID>2285 </input>
<output>
<ID>OUT_0</ID>2291 </output>
<input>
<ID>clear</ID>2246 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1998</ID>
<type>AE_SMALL_INVERTER</type>
<position>-841.5,-4078</position>
<input>
<ID>IN_0</ID>2286 </input>
<output>
<ID>OUT_0</ID>2292 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1999</ID>
<type>AE_SMALL_INVERTER</type>
<position>-826.5,-4078</position>
<input>
<ID>IN_0</ID>2287 </input>
<output>
<ID>OUT_0</ID>2293 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2000</ID>
<type>AE_SMALL_INVERTER</type>
<position>-811.5,-4078</position>
<input>
<ID>IN_0</ID>2288 </input>
<output>
<ID>OUT_0</ID>2294 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2001</ID>
<type>AE_SMALL_INVERTER</type>
<position>-800,-4077.5</position>
<input>
<ID>IN_0</ID>2289 </input>
<output>
<ID>OUT_0</ID>2295 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2002</ID>
<type>AE_SMALL_INVERTER</type>
<position>-787,-4078</position>
<input>
<ID>IN_0</ID>2290 </input>
<output>
<ID>OUT_0</ID>2296 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2003</ID>
<type>AE_SMALL_INVERTER</type>
<position>-774,-4077.5</position>
<input>
<ID>IN_0</ID>2291 </input>
<output>
<ID>OUT_0</ID>2297 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2004</ID>
<type>AA_AND4</type>
<position>-823.5,-4094.5</position>
<input>
<ID>IN_0</ID>2295 </input>
<input>
<ID>IN_1</ID>2294 </input>
<input>
<ID>IN_2</ID>2293 </input>
<input>
<ID>IN_3</ID>2292 </input>
<output>
<ID>OUT</ID>2298 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2005</ID>
<type>AA_LABEL</type>
<position>-933,-3964</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2006</ID>
<type>AA_AND2</type>
<position>-787,-4093.5</position>
<input>
<ID>IN_0</ID>2297 </input>
<input>
<ID>IN_1</ID>2296 </input>
<output>
<ID>OUT</ID>2303 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2007</ID>
<type>AA_AND2</type>
<position>-809.5,-4116.5</position>
<input>
<ID>IN_0</ID>2303 </input>
<input>
<ID>IN_1</ID>2298 </input>
<output>
<ID>OUT</ID>2244 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2008</ID>
<type>AI_XOR2</type>
<position>-852.5,-4061.5</position>
<input>
<ID>IN_0</ID>2203 </input>
<input>
<ID>IN_1</ID>2336 </input>
<output>
<ID>OUT</ID>2280 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2009</ID>
<type>AI_XOR2</type>
<position>-839,-4061.5</position>
<input>
<ID>IN_0</ID>2207 </input>
<input>
<ID>IN_1</ID>2338 </input>
<output>
<ID>OUT</ID>2281 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2010</ID>
<type>AI_XOR2</type>
<position>-826,-4061.5</position>
<input>
<ID>IN_0</ID>2220 </input>
<input>
<ID>IN_1</ID>2340 </input>
<output>
<ID>OUT</ID>2282 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2011</ID>
<type>AI_XOR2</type>
<position>-813,-4061.5</position>
<input>
<ID>IN_0</ID>2223 </input>
<input>
<ID>IN_1</ID>2342 </input>
<output>
<ID>OUT</ID>2283 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2012</ID>
<type>AI_XOR2</type>
<position>-800.5,-4062</position>
<input>
<ID>IN_0</ID>2228 </input>
<input>
<ID>IN_1</ID>2344 </input>
<output>
<ID>OUT</ID>2284 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2013</ID>
<type>AA_AND2</type>
<position>-763.5,-4452.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2277 </input>
<output>
<ID>OUT</ID>2300 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2014</ID>
<type>AI_XOR2</type>
<position>-788,-4062</position>
<input>
<ID>IN_0</ID>2229 </input>
<input>
<ID>IN_1</ID>2346 </input>
<output>
<ID>OUT</ID>2285 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2015</ID>
<type>AA_LABEL</type>
<position>-991.5,-3938</position>
<gparam>LABEL_TEXT Zone 4</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2016</ID>
<type>AA_AND2</type>
<position>-762.5,-4443</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2277 </input>
<output>
<ID>OUT</ID>2301 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2017</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-873.5,-4024.5</position>
<input>
<ID>J</ID>2327 </input>
<output>
<ID>Q</ID>2336 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2347 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2018</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-886.5,-4014.5</position>
<input>
<ID>J</ID>2337 </input>
<output>
<ID>Q</ID>2338 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2347 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2019</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-899.5,-4003.5</position>
<input>
<ID>J</ID>2339 </input>
<output>
<ID>Q</ID>2340 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2347 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2020</ID>
<type>AI_XOR2</type>
<position>-796,-4109.5</position>
<input>
<ID>IN_0</ID>2298 </input>
<input>
<ID>IN_1</ID>2303 </input>
<output>
<ID>OUT</ID>2162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2021</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-907,-3994.5</position>
<input>
<ID>J</ID>2341 </input>
<output>
<ID>Q</ID>2342 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2347 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2022</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-915.5,-3987</position>
<input>
<ID>J</ID>2343 </input>
<output>
<ID>Q</ID>2344 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2347 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2023</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-924.5,-3979.5</position>
<input>
<ID>J</ID>2345 </input>
<output>
<ID>Q</ID>2346 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2347 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2024</ID>
<type>CC_PULSE</type>
<position>-933,-3971.5</position>
<output>
<ID>OUT_0</ID>2347 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2025</ID>
<type>AA_AND2</type>
<position>-938.5,-4022.5</position>
<input>
<ID>IN_0</ID>2279 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2327 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2026</ID>
<type>AA_AND2</type>
<position>-939,-4012.5</position>
<input>
<ID>IN_0</ID>2279 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2027</ID>
<type>AA_AND2</type>
<position>-940.5,-4001.5</position>
<input>
<ID>IN_0</ID>2279 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2339 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2028</ID>
<type>AA_AND2</type>
<position>-941,-3992.5</position>
<input>
<ID>IN_0</ID>2279 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2029</ID>
<type>AA_AND2</type>
<position>-762,-4434.5</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2277 </input>
<output>
<ID>OUT</ID>2302 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2030</ID>
<type>AA_AND2</type>
<position>-761,-4426</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2277 </input>
<output>
<ID>OUT</ID>2304 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2031</ID>
<type>AI_XOR2</type>
<position>-767,-4532.5</position>
<input>
<ID>IN_0</ID>2305 </input>
<input>
<ID>IN_1</ID>2306 </input>
<output>
<ID>OUT</ID>2307 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2032</ID>
<type>AI_XOR2</type>
<position>-1354.5,-3191</position>
<input>
<ID>IN_0</ID>2328 </input>
<input>
<ID>IN_1</ID>2662 </input>
<output>
<ID>OUT</ID>2666 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2033</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-792,-4550</position>
<input>
<ID>J</ID>2306 </input>
<output>
<ID>Q</ID>2308 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2034</ID>
<type>AA_AND2</type>
<position>-778,-4551.5</position>
<input>
<ID>IN_0</ID>2308 </input>
<input>
<ID>IN_1</ID>2572 </input>
<output>
<ID>OUT</ID>2310 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2035</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-891.5,-3618.5</position>
<input>
<ID>J</ID>2664 </input>
<output>
<ID>Q</ID>2661 </output>
<input>
<ID>clear</ID>2664 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2665 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2036</ID>
<type>AA_AND2</type>
<position>-774,-4707.5</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2310 </input>
<output>
<ID>OUT</ID>2309 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2037</ID>
<type>AA_AND2</type>
<position>-952,-3635</position>
<input>
<ID>IN_0</ID>2415 </input>
<input>
<ID>IN_1</ID>2668 </input>
<output>
<ID>OUT</ID>2663 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2038</ID>
<type>AA_AND2</type>
<position>-763,-4698</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2310 </input>
<output>
<ID>OUT</ID>2311 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2039</ID>
<type>AA_AND2</type>
<position>-942,-3985</position>
<input>
<ID>IN_0</ID>2279 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2343 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2040</ID>
<type>AA_AND2</type>
<position>-763.5,-4688.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2310 </input>
<output>
<ID>OUT</ID>2660 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2041</ID>
<type>AE_SMALL_INVERTER</type>
<position>-909.5,-3624.5</position>
<input>
<ID>IN_0</ID>2663 </input>
<output>
<ID>OUT_0</ID>2664 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2042</ID>
<type>AA_AND2</type>
<position>-763,-4680</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2310 </input>
<output>
<ID>OUT</ID>2312 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2043</ID>
<type>GA_LED</type>
<position>-884.5,-3620.5</position>
<input>
<ID>N_in0</ID>2665 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2044</ID>
<type>AA_AND2</type>
<position>-763,-4671.5</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2310 </input>
<output>
<ID>OUT</ID>2313 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2045</ID>
<type>AA_TOGGLE</type>
<position>-917.5,-3475</position>
<output>
<ID>OUT_0</ID>2667 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2046</ID>
<type>AA_AND2</type>
<position>-762.5,-4664</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2310 </input>
<output>
<ID>OUT</ID>2314 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2047</ID>
<type>AA_AND2</type>
<position>-941,-3631</position>
<input>
<ID>IN_0</ID>2414 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2668 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2048</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-894.5,-3743</position>
<input>
<ID>J</ID>2670 </input>
<output>
<ID>Q</ID>2673 </output>
<input>
<ID>clear</ID>2670 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2671 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2049</ID>
<type>AA_AND2</type>
<position>-964.5,-3754</position>
<input>
<ID>IN_0</ID>2386 </input>
<input>
<ID>IN_1</ID>2672 </input>
<output>
<ID>OUT</ID>2669 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2050</ID>
<type>AE_SMALL_INVERTER</type>
<position>-971.5,-3752</position>
<input>
<ID>IN_0</ID>2669 </input>
<output>
<ID>OUT_0</ID>2670 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2051</ID>
<type>BA_NAND2</type>
<position>-580.5,-3633.5</position>
<input>
<ID>IN_0</ID>2307 </input>
<input>
<ID>IN_1</ID>2306 </input>
<output>
<ID>OUT</ID>2331 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2052</ID>
<type>GA_LED</type>
<position>-887.5,-3745</position>
<input>
<ID>N_in0</ID>2671 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2053</ID>
<type>AI_XOR2</type>
<position>-765.5,-4765.5</position>
<input>
<ID>IN_0</ID>2315 </input>
<input>
<ID>IN_1</ID>2316 </input>
<output>
<ID>OUT</ID>2317 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2054</ID>
<type>AA_AND2</type>
<position>-952.5,-3753</position>
<input>
<ID>IN_0</ID>2385 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2672 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2055</ID>
<type>BA_NAND2</type>
<position>-567.5,-3633.5</position>
<input>
<ID>IN_0</ID>2317 </input>
<input>
<ID>IN_1</ID>2316 </input>
<output>
<ID>OUT</ID>2332 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2056</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-787.5,-4784.5</position>
<input>
<ID>J</ID>2316 </input>
<output>
<ID>Q</ID>2318 </output>
<input>
<ID>clear</ID>2667 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2057</ID>
<type>AA_AND2</type>
<position>-772,-4789</position>
<input>
<ID>IN_0</ID>2318 </input>
<input>
<ID>IN_1</ID>2606 </input>
<output>
<ID>OUT</ID>2320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2058</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-918.5,-3914</position>
<input>
<ID>J</ID>2675 </input>
<output>
<ID>Q</ID>2678 </output>
<input>
<ID>clear</ID>2675 </input>
<input>
<ID>clock</ID>2486 </input>
<output>
<ID>nQ</ID>2676 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2059</ID>
<type>AA_AND2</type>
<position>-756.5,-4929</position>
<input>
<ID>IN_0</ID>2530 </input>
<input>
<ID>IN_1</ID>2320 </input>
<output>
<ID>OUT</ID>2319 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2060</ID>
<type>AA_AND2</type>
<position>-929,-3924</position>
<input>
<ID>IN_0</ID>2227 </input>
<input>
<ID>IN_1</ID>2677 </input>
<output>
<ID>OUT</ID>2674 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2061</ID>
<type>AE_SMALL_INVERTER</type>
<position>-936.5,-3920</position>
<input>
<ID>IN_0</ID>2674 </input>
<output>
<ID>OUT_0</ID>2675 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2062</ID>
<type>AA_AND2</type>
<position>-744.5,-4920.5</position>
<input>
<ID>IN_0</ID>2531 </input>
<input>
<ID>IN_1</ID>2320 </input>
<output>
<ID>OUT</ID>2321 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2063</ID>
<type>GA_LED</type>
<position>-911.5,-3916</position>
<input>
<ID>N_in0</ID>2676 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2064</ID>
<type>AA_AND2</type>
<position>-743,-4910.5</position>
<input>
<ID>IN_0</ID>2532 </input>
<input>
<ID>IN_1</ID>2320 </input>
<output>
<ID>OUT</ID>2322 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2065</ID>
<type>AA_AND2</type>
<position>-888.5,-3922</position>
<input>
<ID>IN_0</ID>2226 </input>
<input>
<ID>IN_1</ID>2667 </input>
<output>
<ID>OUT</ID>2677 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2066</ID>
<type>AA_TOGGLE</type>
<position>-982.5,-3490</position>
<output>
<ID>OUT_0</ID>2690 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2067</ID>
<type>AA_AND2</type>
<position>-943,-3977.5</position>
<input>
<ID>IN_0</ID>2279 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2068</ID>
<type>AA_LABEL</type>
<position>-979,-3485</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2069</ID>
<type>AE_DFF_LOW</type>
<position>-848.5,-4070</position>
<input>
<ID>IN_0</ID>2280 </input>
<output>
<ID>OUT_0</ID>2286 </output>
<input>
<ID>clear</ID>2246 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2070</ID>
<type>AE_DFF_LOW</type>
<position>-822,-4269.5</position>
<input>
<ID>IN_0</ID>2351 </input>
<output>
<ID>OUT_0</ID>2357 </output>
<input>
<ID>clear</ID>2251 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2071</ID>
<type>AI_XOR2</type>
<position>-990,-3500</position>
<input>
<ID>IN_0</ID>2690 </input>
<input>
<ID>IN_1</ID>2689 </input>
<output>
<ID>OUT</ID>2393 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2072</ID>
<type>AE_DFF_LOW</type>
<position>-808.5,-4269.5</position>
<input>
<ID>IN_0</ID>2352 </input>
<output>
<ID>OUT_0</ID>2358 </output>
<input>
<ID>clear</ID>2251 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2073</ID>
<type>AE_DFF_LOW</type>
<position>-793.5,-4269.5</position>
<input>
<ID>IN_0</ID>2353 </input>
<output>
<ID>OUT_0</ID>2359 </output>
<input>
<ID>clear</ID>2251 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2074</ID>
<type>AI_XOR2</type>
<position>-985,-3652</position>
<input>
<ID>IN_0</ID>2692 </input>
<input>
<ID>IN_1</ID>2691 </input>
<output>
<ID>OUT</ID>2544 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2075</ID>
<type>AE_DFF_LOW</type>
<position>-783,-4269.5</position>
<input>
<ID>IN_0</ID>2354 </input>
<output>
<ID>OUT_0</ID>2360 </output>
<input>
<ID>clear</ID>2251 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2076</ID>
<type>AE_DFF_LOW</type>
<position>-770,-4269.5</position>
<input>
<ID>IN_0</ID>2355 </input>
<output>
<ID>OUT_0</ID>2361 </output>
<input>
<ID>clear</ID>2251 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2077</ID>
<type>AA_TOGGLE</type>
<position>-983.5,-3643.5</position>
<output>
<ID>OUT_0</ID>2692 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2078</ID>
<type>AE_SMALL_INVERTER</type>
<position>-831,-4277</position>
<input>
<ID>IN_0</ID>2356 </input>
<output>
<ID>OUT_0</ID>2362 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2079</ID>
<type>AE_SMALL_INVERTER</type>
<position>-816,-4277</position>
<input>
<ID>IN_0</ID>2357 </input>
<output>
<ID>OUT_0</ID>2363 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2080</ID>
<type>AA_LABEL</type>
<position>-982.5,-3639.5</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2081</ID>
<type>AE_SMALL_INVERTER</type>
<position>-801,-4277</position>
<input>
<ID>IN_0</ID>2358 </input>
<output>
<ID>OUT_0</ID>2364 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2082</ID>
<type>AI_XOR2</type>
<position>-994,-3775.5</position>
<input>
<ID>IN_0</ID>2694 </input>
<input>
<ID>IN_1</ID>2693 </input>
<output>
<ID>OUT</ID>2174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2083</ID>
<type>AE_SMALL_INVERTER</type>
<position>-789.5,-4276.5</position>
<input>
<ID>IN_0</ID>2359 </input>
<output>
<ID>OUT_0</ID>2365 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2084</ID>
<type>AA_TOGGLE</type>
<position>-992.5,-3767</position>
<output>
<ID>OUT_0</ID>2694 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2085</ID>
<type>AE_SMALL_INVERTER</type>
<position>-776.5,-4277</position>
<input>
<ID>IN_0</ID>2360 </input>
<output>
<ID>OUT_0</ID>2366 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2086</ID>
<type>AA_LABEL</type>
<position>-991.5,-3763</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2087</ID>
<type>AE_SMALL_INVERTER</type>
<position>-763.5,-4276.5</position>
<input>
<ID>IN_0</ID>2361 </input>
<output>
<ID>OUT_0</ID>2367 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2088</ID>
<type>AA_TOGGLE</type>
<position>-999,-3767</position>
<output>
<ID>OUT_0</ID>2693 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2089</ID>
<type>AI_XOR2</type>
<position>-980.5,-3952</position>
<input>
<ID>IN_0</ID>2696 </input>
<input>
<ID>IN_1</ID>2695 </input>
<output>
<ID>OUT</ID>2279 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2091</ID>
<type>AA_AND4</type>
<position>-813,-4293.5</position>
<input>
<ID>IN_0</ID>2365 </input>
<input>
<ID>IN_1</ID>2364 </input>
<input>
<ID>IN_2</ID>2363 </input>
<input>
<ID>IN_3</ID>2362 </input>
<output>
<ID>OUT</ID>2368 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2093</ID>
<type>AA_TOGGLE</type>
<position>-977.5,-3943</position>
<output>
<ID>OUT_0</ID>2696 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2095</ID>
<type>AA_LABEL</type>
<position>-922.5,-4163</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2097</ID>
<type>AA_LABEL</type>
<position>-971.5,-3939</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2099</ID>
<type>AA_AND2</type>
<position>-776.5,-4292.5</position>
<input>
<ID>IN_0</ID>2367 </input>
<input>
<ID>IN_1</ID>2366 </input>
<output>
<ID>OUT</ID>2369 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2101</ID>
<type>AA_TOGGLE</type>
<position>-984.5,-3943</position>
<output>
<ID>OUT_0</ID>2695 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2103</ID>
<type>AA_AND2</type>
<position>-799,-4315.5</position>
<input>
<ID>IN_0</ID>2369 </input>
<input>
<ID>IN_1</ID>2368 </input>
<output>
<ID>OUT</ID>2274 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2105</ID>
<type>AI_XOR2</type>
<position>-961,-4149</position>
<input>
<ID>IN_0</ID>2698 </input>
<input>
<ID>IN_1</ID>2697 </input>
<output>
<ID>OUT</ID>2349 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2107</ID>
<type>AI_XOR2</type>
<position>-842,-4260.5</position>
<input>
<ID>IN_0</ID>2266 </input>
<input>
<ID>IN_1</ID>2371 </input>
<output>
<ID>OUT</ID>2350 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2109</ID>
<type>AA_TOGGLE</type>
<position>-959.5,-4140.5</position>
<output>
<ID>OUT_0</ID>2698 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2110</ID>
<type>AI_XOR2</type>
<position>-828.5,-4260.5</position>
<input>
<ID>IN_0</ID>2268 </input>
<input>
<ID>IN_1</ID>2373 </input>
<output>
<ID>OUT</ID>2351 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2111</ID>
<type>AA_LABEL</type>
<position>-958.5,-4136.5</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2112</ID>
<type>AI_XOR2</type>
<position>-815.5,-4260.5</position>
<input>
<ID>IN_0</ID>2269 </input>
<input>
<ID>IN_1</ID>2375 </input>
<output>
<ID>OUT</ID>2352 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2113</ID>
<type>AA_TOGGLE</type>
<position>-966,-4140.5</position>
<output>
<ID>OUT_0</ID>2697 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2114</ID>
<type>AI_XOR2</type>
<position>-802.5,-4260.5</position>
<input>
<ID>IN_0</ID>2270 </input>
<input>
<ID>IN_1</ID>2377 </input>
<output>
<ID>OUT</ID>2353 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2115</ID>
<type>AI_XOR2</type>
<position>-967.5,-4366.5</position>
<input>
<ID>IN_0</ID>2700 </input>
<input>
<ID>IN_1</ID>2699 </input>
<output>
<ID>OUT</ID>2387 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2116</ID>
<type>AI_XOR2</type>
<position>-790,-4261</position>
<input>
<ID>IN_0</ID>2271 </input>
<input>
<ID>IN_1</ID>2379 </input>
<output>
<ID>OUT</ID>2354 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2117</ID>
<type>AA_TOGGLE</type>
<position>-966,-4358</position>
<output>
<ID>OUT_0</ID>2700 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2118</ID>
<type>AA_AND2</type>
<position>-742.5,-4901</position>
<input>
<ID>IN_0</ID>2533 </input>
<input>
<ID>IN_1</ID>2320 </input>
<output>
<ID>OUT</ID>2323 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2119</ID>
<type>AA_LABEL</type>
<position>-965,-4354</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2120</ID>
<type>AI_XOR2</type>
<position>-777.5,-4261</position>
<input>
<ID>IN_0</ID>2272 </input>
<input>
<ID>IN_1</ID>2381 </input>
<output>
<ID>OUT</ID>2355 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2121</ID>
<type>AA_TOGGLE</type>
<position>-972.5,-4358</position>
<output>
<ID>OUT_0</ID>2699 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2122</ID>
<type>AI_XOR2</type>
<position>-966.5,-4608.5</position>
<input>
<ID>IN_0</ID>2702 </input>
<input>
<ID>IN_1</ID>2701 </input>
<output>
<ID>OUT</ID>2572 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2123</ID>
<type>AA_LABEL</type>
<position>-973,-4132.5</position>
<gparam>LABEL_TEXT Zone 5</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2124</ID>
<type>AA_TOGGLE</type>
<position>-965,-4600</position>
<output>
<ID>OUT_0</ID>2702 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2125</ID>
<type>AA_AND2</type>
<position>-743,-4892.5</position>
<input>
<ID>IN_0</ID>2534 </input>
<input>
<ID>IN_1</ID>2320 </input>
<output>
<ID>OUT</ID>2324 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2126</ID>
<type>AA_LABEL</type>
<position>-964,-4596</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2127</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-863,-4223.5</position>
<input>
<ID>J</ID>2370 </input>
<output>
<ID>Q</ID>2371 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2382 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2128</ID>
<type>AA_TOGGLE</type>
<position>-971.5,-4600</position>
<output>
<ID>OUT_0</ID>2701 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2129</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-876,-4213.5</position>
<input>
<ID>J</ID>2372 </input>
<output>
<ID>Q</ID>2373 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2382 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2130</ID>
<type>AI_XOR2</type>
<position>-959.5,-4822</position>
<input>
<ID>IN_0</ID>2704 </input>
<input>
<ID>IN_1</ID>2703 </input>
<output>
<ID>OUT</ID>2606 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2131</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-889,-4202.5</position>
<input>
<ID>J</ID>2374 </input>
<output>
<ID>Q</ID>2375 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2382 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2132</ID>
<type>AA_TOGGLE</type>
<position>-958,-4813.5</position>
<output>
<ID>OUT_0</ID>2704 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2133</ID>
<type>AI_XOR2</type>
<position>-785.5,-4308.5</position>
<input>
<ID>IN_0</ID>2368 </input>
<input>
<ID>IN_1</ID>2369 </input>
<output>
<ID>OUT</ID>2164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2134</ID>
<type>AA_LABEL</type>
<position>-957,-4809.5</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2135</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-896.5,-4193.5</position>
<input>
<ID>J</ID>2376 </input>
<output>
<ID>Q</ID>2377 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2382 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2136</ID>
<type>AA_TOGGLE</type>
<position>-964.5,-4813.5</position>
<output>
<ID>OUT_0</ID>2703 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2137</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-905,-4186</position>
<input>
<ID>J</ID>2378 </input>
<output>
<ID>Q</ID>2379 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2382 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2138</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-914,-4178.5</position>
<input>
<ID>J</ID>2380 </input>
<output>
<ID>Q</ID>2381 </output>
<input>
<ID>clear</ID>2653 </input>
<input>
<ID>clock</ID>2382 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2139</ID>
<type>GA_LED</type>
<position>-959.5,-3490</position>
<input>
<ID>N_in0</ID>2690 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2140</ID>
<type>CC_PULSE</type>
<position>-922,-4170.5</position>
<output>
<ID>OUT_0</ID>2382 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2141</ID>
<type>AA_AND2</type>
<position>-928,-4221.5</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2142</ID>
<type>GA_LED</type>
<position>-971.5,-3644.5</position>
<input>
<ID>N_in0</ID>2692 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2143</ID>
<type>AA_AND2</type>
<position>-928.5,-4211.5</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2372 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2144</ID>
<type>GA_LED</type>
<position>-981,-3767.5</position>
<input>
<ID>N_in0</ID>2694 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2145</ID>
<type>AA_AND2</type>
<position>-930,-4200.5</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2146</ID>
<type>GA_LED</type>
<position>-965,-3945</position>
<input>
<ID>N_in0</ID>2696 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2147</ID>
<type>AA_AND2</type>
<position>-930.5,-4191.5</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2376 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2148</ID>
<type>GA_LED</type>
<position>-948,-4143</position>
<input>
<ID>N_in0</ID>2698 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2149</ID>
<type>AA_AND2</type>
<position>-931.5,-4184</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2378 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2150</ID>
<type>GA_LED</type>
<position>-955.5,-4361.5</position>
<input>
<ID>N_in0</ID>2700 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2151</ID>
<type>AA_AND2</type>
<position>-932.5,-4176.5</position>
<input>
<ID>IN_0</ID>2349 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2152</ID>
<type>GA_LED</type>
<position>-954,-4602.5</position>
<input>
<ID>N_in0</ID>2702 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2153</ID>
<type>AE_DFF_LOW</type>
<position>-838,-4269</position>
<input>
<ID>IN_0</ID>2350 </input>
<output>
<ID>OUT_0</ID>2356 </output>
<input>
<ID>clear</ID>2251 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2154</ID>
<type>GA_LED</type>
<position>-948,-4816.5</position>
<input>
<ID>N_in0</ID>2704 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2155</ID>
<type>AE_DFF_LOW</type>
<position>-828.5,-4491.5</position>
<input>
<ID>IN_0</ID>2389 </input>
<output>
<ID>OUT_0</ID>2416 </output>
<input>
<ID>clear</ID>2256 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2156</ID>
<type>AE_DFF_LOW</type>
<position>-814.5,-4491.5</position>
<input>
<ID>IN_0</ID>2390 </input>
<output>
<ID>OUT_0</ID>2417 </output>
<input>
<ID>clear</ID>2256 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2157</ID>
<type>AE_DFF_LOW</type>
<position>-800,-4491.5</position>
<input>
<ID>IN_0</ID>2391 </input>
<output>
<ID>OUT_0</ID>2418 </output>
<input>
<ID>clear</ID>2256 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2158</ID>
<type>AE_DFF_LOW</type>
<position>-789.5,-4491.5</position>
<input>
<ID>IN_0</ID>2392 </input>
<output>
<ID>OUT_0</ID>2489 </output>
<input>
<ID>clear</ID>2256 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2159</ID>
<type>AA_AND4</type>
<position>-841.5,-3750.5</position>
<input>
<ID>IN_0</ID>2200 </input>
<input>
<ID>IN_1</ID>2199 </input>
<input>
<ID>IN_2</ID>2198 </input>
<input>
<ID>IN_3</ID>2197 </input>
<output>
<ID>OUT</ID>2385 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2160</ID>
<type>AA_AND2</type>
<position>-805,-3749.5</position>
<input>
<ID>IN_0</ID>2384 </input>
<input>
<ID>IN_1</ID>2383 </input>
<output>
<ID>OUT</ID>2386 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2161</ID>
<type>AA_AND2</type>
<position>-826,-3767.5</position>
<input>
<ID>IN_0</ID>2386 </input>
<input>
<ID>IN_1</ID>2385 </input>
<output>
<ID>OUT</ID>2687 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2162</ID>
<type>AI_XOR2</type>
<position>-870.5,-3717.5</position>
<input>
<ID>IN_0</ID>2680 </input>
<input>
<ID>IN_1</ID>2640 </input>
<output>
<ID>OUT</ID>2185 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2163</ID>
<type>AI_XOR2</type>
<position>-857,-3717.5</position>
<input>
<ID>IN_0</ID>2681 </input>
<input>
<ID>IN_1</ID>2642 </input>
<output>
<ID>OUT</ID>2186 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2164</ID>
<type>AI_XOR2</type>
<position>-844,-3717.5</position>
<input>
<ID>IN_0</ID>2682 </input>
<input>
<ID>IN_1</ID>2644 </input>
<output>
<ID>OUT</ID>2187 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2165</ID>
<type>AI_XOR2</type>
<position>-831,-3717.5</position>
<input>
<ID>IN_0</ID>2683 </input>
<input>
<ID>IN_1</ID>2646 </input>
<output>
<ID>OUT</ID>2188 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2166</ID>
<type>AI_XOR2</type>
<position>-818.5,-3718</position>
<input>
<ID>IN_0</ID>2684 </input>
<input>
<ID>IN_1</ID>2648 </input>
<output>
<ID>OUT</ID>2189 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2167</ID>
<type>AI_XOR2</type>
<position>-806,-3718</position>
<input>
<ID>IN_0</ID>2685 </input>
<input>
<ID>IN_1</ID>2650 </input>
<output>
<ID>OUT</ID>2190 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2168</ID>
<type>AE_DFF_LOW</type>
<position>-866.5,-3726</position>
<input>
<ID>IN_0</ID>2185 </input>
<output>
<ID>OUT_0</ID>2191 </output>
<input>
<ID>clear</ID>2673 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2169</ID>
<type>AE_DFF_LOW</type>
<position>-776.5,-4491.5</position>
<input>
<ID>IN_0</ID>2394 </input>
<output>
<ID>OUT_0</ID>2496 </output>
<input>
<ID>clear</ID>2256 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2170</ID>
<type>AE_SMALL_INVERTER</type>
<position>-837.5,-4499</position>
<input>
<ID>IN_0</ID>2395 </input>
<output>
<ID>OUT_0</ID>2497 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2171</ID>
<type>AA_AND2</type>
<position>-956,-3553.5</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2433 </input>
<output>
<ID>OUT</ID>2552 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2172</ID>
<type>AE_SMALL_INVERTER</type>
<position>-822.5,-4499</position>
<input>
<ID>IN_0</ID>2416 </input>
<output>
<ID>OUT_0</ID>2538 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2173</ID>
<type>AE_SMALL_INVERTER</type>
<position>-807.5,-4499</position>
<input>
<ID>IN_0</ID>2417 </input>
<output>
<ID>OUT_0</ID>2539 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2174</ID>
<type>AA_AND2</type>
<position>-956.5,-3543.5</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2451 </input>
<output>
<ID>OUT</ID>2554 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2175</ID>
<type>AA_AND2</type>
<position>-958,-3532.5</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2452 </input>
<output>
<ID>OUT</ID>2556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2176</ID>
<type>AE_SMALL_INVERTER</type>
<position>-796,-4498.5</position>
<input>
<ID>IN_0</ID>2418 </input>
<output>
<ID>OUT_0</ID>2540 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2177</ID>
<type>AA_AND2</type>
<position>-958.5,-3523.5</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2453 </input>
<output>
<ID>OUT</ID>2558 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2178</ID>
<type>AE_SMALL_INVERTER</type>
<position>-783,-4499</position>
<input>
<ID>IN_0</ID>2489 </input>
<output>
<ID>OUT_0</ID>2541 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2179</ID>
<type>AE_SMALL_INVERTER</type>
<position>-770,-4498.5</position>
<input>
<ID>IN_0</ID>2496 </input>
<output>
<ID>OUT_0</ID>2542 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2180</ID>
<type>AA_AND2</type>
<position>-959.5,-3516</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2454 </input>
<output>
<ID>OUT</ID>2560 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2181</ID>
<type>AA_AND2</type>
<position>-960.5,-3508.5</position>
<input>
<ID>IN_0</ID>2393 </input>
<input>
<ID>IN_1</ID>2455 </input>
<output>
<ID>OUT</ID>2562 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2182</ID>
<type>AA_LABEL</type>
<position>-1247,-3511.5</position>
<gparam>LABEL_TEXT Checking condition for 60</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2183</ID>
<type>AA_TOGGLE</type>
<position>-1377.5,-3372.5</position>
<output>
<ID>OUT_0</ID>2420 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2184</ID>
<type>AA_LABEL</type>
<position>-1045.5,-3430.5</position>
<gparam>LABEL_TEXT Problematic Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2185</ID>
<type>BA_NAND4</type>
<position>-1068.5,-3375.5</position>
<input>
<ID>IN_0</ID>2437 </input>
<input>
<ID>IN_1</ID>2441 </input>
<input>
<ID>IN_2</ID>2445 </input>
<input>
<ID>IN_3</ID>2450 </input>
<output>
<ID>OUT</ID>2427 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2186</ID>
<type>AE_DFF_LOW</type>
<position>-1267.5,-3445.5</position>
<input>
<ID>IN_0</ID>2428 </input>
<output>
<ID>OUT_0</ID>2433 </output>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2187</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1285.5,-3401</position>
<input>
<ID>J</ID>2456 </input>
<input>
<ID>K</ID>2458 </input>
<output>
<ID>Q</ID>2428 </output>
<input>
<ID>clear</ID>2427 </input>
<input>
<ID>clock</ID>2449 </input>
<output>
<ID>nQ</ID>2429 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2188</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1236,-3401.5</position>
<input>
<ID>J</ID>2468 </input>
<input>
<ID>K</ID>2469 </input>
<output>
<ID>Q</ID>2432 </output>
<input>
<ID>clear</ID>2427 </input>
<input>
<ID>clock</ID>2449 </input>
<output>
<ID>nQ</ID>2435 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2189</ID>
<type>AE_DFF_LOW</type>
<position>-1224.5,-3445</position>
<input>
<ID>IN_0</ID>2432 </input>
<output>
<ID>OUT_0</ID>2451 </output>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2190</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1210,-3401</position>
<input>
<ID>J</ID>2470 </input>
<input>
<ID>K</ID>2471 </input>
<output>
<ID>Q</ID>2437 </output>
<input>
<ID>clear</ID>2427 </input>
<input>
<ID>clock</ID>2449 </input>
<output>
<ID>nQ</ID>2440 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2191</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1180,-3401.5</position>
<input>
<ID>J</ID>2472 </input>
<input>
<ID>K</ID>2473 </input>
<output>
<ID>Q</ID>2441 </output>
<input>
<ID>clear</ID>2427 </input>
<input>
<ID>clock</ID>2449 </input>
<output>
<ID>nQ</ID>2442 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2192</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1141.5,-3403.5</position>
<input>
<ID>J</ID>2474 </input>
<input>
<ID>K</ID>2475 </input>
<output>
<ID>Q</ID>2445 </output>
<input>
<ID>clear</ID>2427 </input>
<input>
<ID>clock</ID>2449 </input>
<output>
<ID>nQ</ID>2446 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2193</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1093,-3404</position>
<input>
<ID>J</ID>2476 </input>
<input>
<ID>K</ID>2477 </input>
<output>
<ID>Q</ID>2450 </output>
<input>
<ID>clear</ID>2427 </input>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2194</ID>
<type>AE_DFF_LOW</type>
<position>-1195,-3445</position>
<input>
<ID>IN_0</ID>2437 </input>
<output>
<ID>OUT_0</ID>2452 </output>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2195</ID>
<type>AA_AND2</type>
<position>-1269,-3392</position>
<input>
<ID>IN_0</ID>2484 </input>
<input>
<ID>IN_1</ID>2428 </input>
<output>
<ID>OUT</ID>2430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2196</ID>
<type>AE_DFF_LOW</type>
<position>-866,-3601</position>
<input>
<ID>IN_0</ID>2396 </input>
<output>
<ID>OUT_0</ID>2402 </output>
<input>
<ID>clear</ID>2661 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2197</ID>
<type>AA_AND2</type>
<position>-1270,-3409.5</position>
<input>
<ID>IN_0</ID>2429 </input>
<input>
<ID>IN_1</ID>2485 </input>
<output>
<ID>OUT</ID>2431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2198</ID>
<type>AA_AND2</type>
<position>-1228,-3392</position>
<input>
<ID>IN_0</ID>2430 </input>
<input>
<ID>IN_1</ID>2432 </input>
<output>
<ID>OUT</ID>2434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2199</ID>
<type>AA_AND2</type>
<position>-1225.5,-3410.5</position>
<input>
<ID>IN_0</ID>2435 </input>
<input>
<ID>IN_1</ID>2431 </input>
<output>
<ID>OUT</ID>2436 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2200</ID>
<type>AA_AND2</type>
<position>-1198.5,-3393.5</position>
<input>
<ID>IN_0</ID>2434 </input>
<input>
<ID>IN_1</ID>2437 </input>
<output>
<ID>OUT</ID>2438 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2201</ID>
<type>AA_AND2</type>
<position>-1196,-3412</position>
<input>
<ID>IN_0</ID>2440 </input>
<input>
<ID>IN_1</ID>2436 </input>
<output>
<ID>OUT</ID>2439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2202</ID>
<type>AA_AND2</type>
<position>-1172,-3394.5</position>
<input>
<ID>IN_0</ID>2438 </input>
<input>
<ID>IN_1</ID>2441 </input>
<output>
<ID>OUT</ID>2443 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2203</ID>
<type>AA_AND2</type>
<position>-1170.5,-3412</position>
<input>
<ID>IN_0</ID>2442 </input>
<input>
<ID>IN_1</ID>2439 </input>
<output>
<ID>OUT</ID>2444 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2204</ID>
<type>AA_AND2</type>
<position>-1125,-3393.5</position>
<input>
<ID>IN_0</ID>2443 </input>
<input>
<ID>IN_1</ID>2445 </input>
<output>
<ID>OUT</ID>2447 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2205</ID>
<type>AA_AND2</type>
<position>-1124.5,-3411</position>
<input>
<ID>IN_0</ID>2446 </input>
<input>
<ID>IN_1</ID>2444 </input>
<output>
<ID>OUT</ID>2448 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2206</ID>
<type>AE_DFF_LOW</type>
<position>-1166.5,-3445</position>
<input>
<ID>IN_0</ID>2441 </input>
<output>
<ID>OUT_0</ID>2453 </output>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2207</ID>
<type>AE_OR2</type>
<position>-1255,-3401.5</position>
<input>
<ID>IN_0</ID>2430 </input>
<input>
<ID>IN_1</ID>2431 </input>
<output>
<ID>OUT</ID>2468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2208</ID>
<type>AE_DFF_LOW</type>
<position>-1120.5,-3445</position>
<input>
<ID>IN_0</ID>2445 </input>
<output>
<ID>OUT_0</ID>2454 </output>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2209</ID>
<type>AE_OR2</type>
<position>-1218.5,-3400.5</position>
<input>
<ID>IN_0</ID>2434 </input>
<input>
<ID>IN_1</ID>2436 </input>
<output>
<ID>OUT</ID>2471 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2210</ID>
<type>AE_OR2</type>
<position>-1190,-3401</position>
<input>
<ID>IN_0</ID>2438 </input>
<input>
<ID>IN_1</ID>2439 </input>
<output>
<ID>OUT</ID>2472 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2211</ID>
<type>AE_OR2</type>
<position>-1161,-3401.5</position>
<input>
<ID>IN_0</ID>2443 </input>
<input>
<ID>IN_1</ID>2444 </input>
<output>
<ID>OUT</ID>2474 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2212</ID>
<type>AE_OR2</type>
<position>-1117,-3402</position>
<input>
<ID>IN_0</ID>2447 </input>
<input>
<ID>IN_1</ID>2448 </input>
<output>
<ID>OUT</ID>2476 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2213</ID>
<type>AE_DFF_LOW</type>
<position>-1072.5,-3445.5</position>
<input>
<ID>IN_0</ID>2450 </input>
<output>
<ID>OUT_0</ID>2455 </output>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2214</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-1068.5,-3425</position>
<input>
<ID>IN_0</ID>2428 </input>
<input>
<ID>IN_1</ID>2432 </input>
<input>
<ID>IN_2</ID>2437 </input>
<input>
<ID>IN_3</ID>2441 </input>
<input>
<ID>IN_4</ID>2445 </input>
<input>
<ID>IN_5</ID>2450 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2215</ID>
<type>AE_DFF_LOW</type>
<position>-1349,-3409.5</position>
<input>
<ID>IN_0</ID>2483 </input>
<output>
<ID>OUTINV_0</ID>2485 </output>
<output>
<ID>OUT_0</ID>2484 </output>
<input>
<ID>clear</ID>2426 </input>
<input>
<ID>clock</ID>2449 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2216</ID>
<type>CC_PULSE</type>
<position>-1396.5,-3404</position>
<output>
<ID>OUT_0</ID>2481 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2217</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-1049,-3455.5</position>
<input>
<ID>IN_0</ID>2433 </input>
<input>
<ID>IN_1</ID>2451 </input>
<input>
<ID>IN_2</ID>2452 </input>
<input>
<ID>IN_3</ID>2453 </input>
<input>
<ID>IN_4</ID>2454 </input>
<input>
<ID>IN_5</ID>2455 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2218</ID>
<type>CC_PULSE</type>
<position>-1395,-3422</position>
<output>
<ID>OUT_0</ID>2480 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2219</ID>
<type>EE_VDD</type>
<position>-1344.5,-3369</position>
<output>
<ID>OUT_0</ID>2479 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2220</ID>
<type>AE_OR2</type>
<position>-1358,-3421</position>
<input>
<ID>IN_0</ID>2481 </input>
<input>
<ID>IN_1</ID>2480 </input>
<output>
<ID>OUT</ID>2449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2221</ID>
<type>AE_DFF_LOW</type>
<position>-850,-3601.5</position>
<input>
<ID>IN_0</ID>2397 </input>
<output>
<ID>OUT_0</ID>2403 </output>
<input>
<ID>clear</ID>2661 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2222</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1375.5,-3404.5</position>
<input>
<ID>IN_0</ID>2481 </input>
<output>
<ID>OUT_0</ID>2482 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2223</ID>
<type>AA_AND2</type>
<position>-1251.5,-3496</position>
<input>
<ID>IN_0</ID>2460 </input>
<input>
<ID>IN_1</ID>2459 </input>
<output>
<ID>OUT</ID>2461 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2224</ID>
<type>AI_XOR2</type>
<position>-1361,-3408.5</position>
<input>
<ID>IN_0</ID>2480 </input>
<input>
<ID>IN_1</ID>2482 </input>
<output>
<ID>OUT</ID>2483 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2225</ID>
<type>AA_LABEL</type>
<position>-1391,-3398</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2226</ID>
<type>AA_AND2</type>
<position>-1177.5,-3482.5</position>
<input>
<ID>IN_0</ID>2462 </input>
<input>
<ID>IN_1</ID>2463 </input>
<output>
<ID>OUT</ID>2464 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2227</ID>
<type>AA_LABEL</type>
<position>-1392,-3427</position>
<gparam>LABEL_TEXT Decrement</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2228</ID>
<type>AA_AND2</type>
<position>-1114.5,-3481</position>
<input>
<ID>IN_0</ID>2465 </input>
<input>
<ID>IN_1</ID>2466 </input>
<output>
<ID>OUT</ID>2467 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2229</ID>
<type>AI_XOR2</type>
<position>-1301,-3390</position>
<input>
<ID>IN_0</ID>2456 </input>
<input>
<ID>IN_1</ID>2457 </input>
<output>
<ID>OUT</ID>2458 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2230</ID>
<type>AE_DFF_LOW</type>
<position>-836.5,-3601.5</position>
<input>
<ID>IN_0</ID>2398 </input>
<output>
<ID>OUT_0</ID>2404 </output>
<input>
<ID>clear</ID>2661 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2231</ID>
<type>AI_XOR2</type>
<position>-1250,-3387.5</position>
<input>
<ID>IN_0</ID>2468 </input>
<input>
<ID>IN_1</ID>2457 </input>
<output>
<ID>OUT</ID>2469 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2232</ID>
<type>AI_XOR2</type>
<position>-1213.5,-3387</position>
<input>
<ID>IN_0</ID>2471 </input>
<input>
<ID>IN_1</ID>2457 </input>
<output>
<ID>OUT</ID>2470 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2233</ID>
<type>AI_XOR2</type>
<position>-1185,-3387.5</position>
<input>
<ID>IN_0</ID>2472 </input>
<input>
<ID>IN_1</ID>2457 </input>
<output>
<ID>OUT</ID>2473 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2234</ID>
<type>AI_XOR2</type>
<position>-1155,-3387.5</position>
<input>
<ID>IN_0</ID>2474 </input>
<input>
<ID>IN_1</ID>2457 </input>
<output>
<ID>OUT</ID>2475 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2235</ID>
<type>AI_XOR2</type>
<position>-1107.5,-3385.5</position>
<input>
<ID>IN_0</ID>2476 </input>
<input>
<ID>IN_1</ID>2457 </input>
<output>
<ID>OUT</ID>2477 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2236</ID>
<type>AA_AND4</type>
<position>-1273,-3518</position>
<input>
<ID>IN_0</ID>2467 </input>
<input>
<ID>IN_1</ID>2464 </input>
<input>
<ID>IN_2</ID>2461 </input>
<input>
<ID>IN_3</ID>2485 </input>
<output>
<ID>OUT</ID>2457 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2237</ID>
<type>AE_DFF_LOW</type>
<position>-821.5,-3601.5</position>
<input>
<ID>IN_0</ID>2399 </input>
<output>
<ID>OUT_0</ID>2405 </output>
<input>
<ID>clear</ID>2661 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2238</ID>
<type>AA_INVERTER</type>
<position>-1257.5,-3473</position>
<input>
<ID>IN_0</ID>2428 </input>
<output>
<ID>OUT_0</ID>2459 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2239</ID>
<type>AA_INVERTER</type>
<position>-1245,-3474</position>
<input>
<ID>IN_0</ID>2432 </input>
<output>
<ID>OUT_0</ID>2460 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2240</ID>
<type>AA_INVERTER</type>
<position>-1181,-3473</position>
<input>
<ID>IN_0</ID>2437 </input>
<output>
<ID>OUT_0</ID>2463 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2241</ID>
<type>AA_INVERTER</type>
<position>-1174,-3473</position>
<input>
<ID>IN_0</ID>2441 </input>
<output>
<ID>OUT_0</ID>2462 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2242</ID>
<type>AE_DFF_LOW</type>
<position>-811,-3601.5</position>
<input>
<ID>IN_0</ID>2400 </input>
<output>
<ID>OUT_0</ID>2406 </output>
<input>
<ID>clear</ID>2661 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2243</ID>
<type>AA_INVERTER</type>
<position>-1116.5,-3472.5</position>
<input>
<ID>IN_0</ID>2445 </input>
<output>
<ID>OUT_0</ID>2466 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2244</ID>
<type>AA_INVERTER</type>
<position>-1111,-3472</position>
<input>
<ID>IN_0</ID>2450 </input>
<output>
<ID>OUT_0</ID>2465 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2245</ID>
<type>AA_LABEL</type>
<position>-1049,-3465.5</position>
<gparam>LABEL_TEXT Actual Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2246</ID>
<type>AA_AND4</type>
<position>-819.5,-4515.5</position>
<input>
<ID>IN_0</ID>2540 </input>
<input>
<ID>IN_1</ID>2539 </input>
<input>
<ID>IN_2</ID>2538 </input>
<input>
<ID>IN_3</ID>2497 </input>
<output>
<ID>OUT</ID>2543 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2247</ID>
<type>AA_AND2</type>
<position>-1351.5,-3375.5</position>
<input>
<ID>IN_0</ID>2479 </input>
<input>
<ID>IN_1</ID>2478 </input>
<output>
<ID>OUT</ID>2456 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2248</ID>
<type>AA_LABEL</type>
<position>-1222.5,-3366</position>
<gparam>LABEL_TEXT Setting Mode</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2249</ID>
<type>AE_DFF_LOW</type>
<position>-798,-3601.5</position>
<input>
<ID>IN_0</ID>2401 </input>
<output>
<ID>OUT_0</ID>2407 </output>
<input>
<ID>clear</ID>2661 </input>
<input>
<ID>clock</ID>2486 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2250</ID>
<type>AA_LABEL</type>
<position>-1357.5,-3362.5</position>
<gparam>LABEL_TEXT On/Off- Settings/Cycle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2251</ID>
<type>AA_LABEL</type>
<position>-929,-4385</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2252</ID>
<type>AA_LABEL</type>
<position>-1390.5,-3182.5</position>
<gparam>LABEL_TEXT Water Button</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2253</ID>
<type>AE_SMALL_INVERTER</type>
<position>-859,-3609</position>
<input>
<ID>IN_0</ID>2402 </input>
<output>
<ID>OUT_0</ID>2408 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2254</ID>
<type>AA_LABEL</type>
<position>-1220.5,-3215</position>
<gparam>LABEL_TEXT Buffer Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2255</ID>
<type>AA_LABEL</type>
<position>-1278.5,-3163.5</position>
<gparam>LABEL_TEXT Seconds Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2256</ID>
<type>AE_SMALL_INVERTER</type>
<position>-844,-3609</position>
<input>
<ID>IN_0</ID>2403 </input>
<output>
<ID>OUT_0</ID>2409 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2257</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1091.5,-3276.5</position>
<input>
<ID>J</ID>2536 </input>
<input>
<ID>K</ID>2657 </input>
<output>
<ID>Q</ID>2487 </output>
<input>
<ID>clear</ID>2348 </input>
<input>
<ID>clock</ID>2508 </input>
<output>
<ID>nQ</ID>2493 </output>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2258</ID>
<type>AA_LABEL</type>
<position>-1222,-3236.5</position>
<gparam>LABEL_TEXT Actual Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2259</ID>
<type>AE_SMALL_INVERTER</type>
<position>-829,-3609</position>
<input>
<ID>IN_0</ID>2404 </input>
<output>
<ID>OUT_0</ID>2410 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2260</ID>
<type>AA_LABEL</type>
<position>-1148,-3255</position>
<gparam>LABEL_TEXT Minutes Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2261</ID>
<type>AE_SMALL_INVERTER</type>
<position>-817.5,-3608.5</position>
<input>
<ID>IN_0</ID>2405 </input>
<output>
<ID>OUT_0</ID>2411 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2262</ID>
<type>AA_LABEL</type>
<position>-1085,-3290.5</position>
<gparam>LABEL_TEXT Buffer Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2263</ID>
<type>AE_SMALL_INVERTER</type>
<position>-804.5,-3609</position>
<input>
<ID>IN_0</ID>2406 </input>
<output>
<ID>OUT_0</ID>2412 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2264</ID>
<type>AI_XOR2</type>
<position>-1206,-3190.5</position>
<input>
<ID>IN_0</ID>2493 </input>
<input>
<ID>IN_1</ID>2495 </input>
<output>
<ID>OUT</ID>2501 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2265</ID>
<type>AA_LABEL</type>
<position>-1201.5,-3180.5</position>
<gparam>LABEL_TEXT Both on seconds counter stop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2266</ID>
<type>AE_SMALL_INVERTER</type>
<position>-791.5,-3608.5</position>
<input>
<ID>IN_0</ID>2407 </input>
<output>
<ID>OUT_0</ID>2413 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2267</ID>
<type>AA_LABEL</type>
<position>-1075.5,-3319.5</position>
<gparam>LABEL_TEXT Actual Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2268</ID>
<type>AI_XOR2</type>
<position>-1107,-3278.5</position>
<input>
<ID>IN_0</ID>2502 </input>
<input>
<ID>IN_1</ID>2487 </input>
<output>
<ID>OUT</ID>2490 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2269</ID>
<type>AA_INVERTER</type>
<position>-1098,-3261.5</position>
<input>
<ID>IN_0</ID>2208 </input>
<output>
<ID>OUT_0</ID>2657 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2270</ID>
<type>AA_AND2</type>
<position>-1344.5,-3214</position>
<input>
<ID>IN_0</ID>2536 </input>
<input>
<ID>IN_1</ID>2486 </input>
<output>
<ID>OUT</ID>2508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2271</ID>
<type>AA_LABEL</type>
<position>-1355.5,-3288</position>
<gparam>LABEL_TEXT Abort</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2272</ID>
<type>AE_OR2</type>
<position>-1291,-3270</position>
<input>
<ID>IN_0</ID>2519 </input>
<input>
<ID>IN_1</ID>2518 </input>
<output>
<ID>OUT</ID>2491 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2273</ID>
<type>AA_TOGGLE</type>
<position>-1357.5,-3284.5</position>
<output>
<ID>OUT_0</ID>2502 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2274</ID>
<type>AE_OR4</type>
<position>-1323,-3261.5</position>
<input>
<ID>IN_0</ID>2517 </input>
<input>
<ID>IN_1</ID>2516 </input>
<input>
<ID>IN_2</ID>2515 </input>
<input>
<ID>IN_3</ID>2514 </input>
<output>
<ID>OUT</ID>2488 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2275</ID>
<type>AE_OR2</type>
<position>-1337,-3267</position>
<input>
<ID>IN_0</ID>2491 </input>
<input>
<ID>IN_1</ID>2488 </input>
<output>
<ID>OUT</ID>2498 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2276</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1332,-3201.5</position>
<input>
<ID>J</ID>2536 </input>
<input>
<ID>K</ID>2536 </input>
<output>
<ID>Q</ID>2507 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2277</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1318.5,-3201.5</position>
<input>
<ID>J</ID>2507 </input>
<input>
<ID>K</ID>2507 </input>
<output>
<ID>Q</ID>2509 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2278</ID>
<type>AA_AND2</type>
<position>-1343.5,-3257.5</position>
<input>
<ID>IN_0</ID>2490 </input>
<input>
<ID>IN_1</ID>2536 </input>
<output>
<ID>OUT</ID>2492 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2279</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1302.5,-3201.5</position>
<input>
<ID>J</ID>2503 </input>
<input>
<ID>K</ID>2503 </input>
<output>
<ID>Q</ID>2511 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2280</ID>
<type>AE_OR2</type>
<position>-1362,-3254.5</position>
<input>
<ID>IN_0</ID>2499 </input>
<input>
<ID>IN_1</ID>2492 </input>
<output>
<ID>OUT</ID>2500 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2281</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1286.5,-3202</position>
<input>
<ID>J</ID>2504 </input>
<input>
<ID>K</ID>2504 </input>
<output>
<ID>Q</ID>2510 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2282</ID>
<type>AA_AND4</type>
<position>-841,-3625.5</position>
<input>
<ID>IN_0</ID>2411 </input>
<input>
<ID>IN_1</ID>2410 </input>
<input>
<ID>IN_2</ID>2409 </input>
<input>
<ID>IN_3</ID>2408 </input>
<output>
<ID>OUT</ID>2414 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2283</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1270.5,-3202.5</position>
<input>
<ID>J</ID>2505 </input>
<input>
<ID>K</ID>2505 </input>
<output>
<ID>Q</ID>2512 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2284</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1253.5,-3202.5</position>
<input>
<ID>J</ID>2506 </input>
<input>
<ID>K</ID>2506 </input>
<output>
<ID>Q</ID>2513 </output>
<input>
<ID>clear</ID>2494 </input>
<input>
<ID>clock</ID>2508 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2285</ID>
<type>AI_XOR2</type>
<position>-1221,-3199.5</position>
<input>
<ID>IN_0</ID>2502 </input>
<input>
<ID>IN_1</ID>2501 </input>
<output>
<ID>OUT</ID>2494 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2286</ID>
<type>AA_TOGGLE</type>
<position>-1369,-3192.5</position>
<output>
<ID>OUT_0</ID>2662 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2287</ID>
<type>AA_LABEL</type>
<position>-1375.5,-3247.5</position>
<gparam>LABEL_TEXT Water On/Off</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2288</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1203.5,-3274.5</position>
<input>
<ID>J</ID>2536 </input>
<input>
<ID>K</ID>2536 </input>
<output>
<ID>Q</ID>2524 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2289</ID>
<type>AA_AND2</type>
<position>-1354.5,-3266</position>
<input>
<ID>IN_0</ID>2498 </input>
<input>
<ID>IN_1</ID>2536 </input>
<output>
<ID>OUT</ID>2499 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2290</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1190,-3274.5</position>
<input>
<ID>J</ID>2524 </input>
<input>
<ID>K</ID>2524 </input>
<output>
<ID>Q</ID>2525 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2291</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-1236,-3216</position>
<input>
<ID>IN_0</ID>2507 </input>
<input>
<ID>IN_1</ID>2509 </input>
<input>
<ID>IN_2</ID>2511 </input>
<input>
<ID>IN_3</ID>2510 </input>
<input>
<ID>IN_4</ID>2512 </input>
<input>
<ID>IN_5</ID>2513 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2292</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1174,-3274.5</position>
<input>
<ID>J</ID>2520 </input>
<input>
<ID>K</ID>2520 </input>
<output>
<ID>Q</ID>2527 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2293</ID>
<type>AA_AND2</type>
<position>-804.5,-3624.5</position>
<input>
<ID>IN_0</ID>2413 </input>
<input>
<ID>IN_1</ID>2412 </input>
<output>
<ID>OUT</ID>2415 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2294</ID>
<type>GA_LED</type>
<position>-1374,-3254.5</position>
<input>
<ID>N_in1</ID>2500 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2295</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1158,-3275</position>
<input>
<ID>J</ID>2521 </input>
<input>
<ID>K</ID>2521 </input>
<output>
<ID>Q</ID>2526 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2296</ID>
<type>AA_AND2</type>
<position>-827,-3647.5</position>
<input>
<ID>IN_0</ID>2415 </input>
<input>
<ID>IN_1</ID>2414 </input>
<output>
<ID>OUT</ID>2655 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2297</ID>
<type>AA_LABEL</type>
<position>-1297.5,-3273.5</position>
<gparam>LABEL_TEXT Conditions for checking whether the counter is running</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2298</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1142,-3274.5</position>
<input>
<ID>J</ID>2522 </input>
<input>
<ID>K</ID>2522 </input>
<output>
<ID>Q</ID>2528 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2299</ID>
<type>BB_CLOCK</type>
<position>-1359,-3215</position>
<output>
<ID>CLK</ID>2486 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 3</lparam></gate>
<gate>
<ID>2300</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-1125,-3274.5</position>
<input>
<ID>J</ID>2523 </input>
<input>
<ID>K</ID>2523 </input>
<output>
<ID>Q</ID>2529 </output>
<input>
<ID>clear</ID>2490 </input>
<input>
<ID>clock</ID>2537 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2301</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-1113,-3289</position>
<input>
<ID>IN_0</ID>2524 </input>
<input>
<ID>IN_1</ID>2525 </input>
<input>
<ID>IN_2</ID>2527 </input>
<input>
<ID>IN_3</ID>2526 </input>
<input>
<ID>IN_4</ID>2528 </input>
<input>
<ID>IN_5</ID>2529 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2302</ID>
<type>AA_AND2</type>
<position>-1311.5,-3191</position>
<input>
<ID>IN_0</ID>2507 </input>
<input>
<ID>IN_1</ID>2509 </input>
<output>
<ID>OUT</ID>2503 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2303</ID>
<type>AA_AND2</type>
<position>-743.5,-4884</position>
<input>
<ID>IN_0</ID>2535 </input>
<input>
<ID>IN_1</ID>2320 </input>
<output>
<ID>OUT</ID>2325 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2304</ID>
<type>AA_AND2</type>
<position>-1183,-3264</position>
<input>
<ID>IN_0</ID>2524 </input>
<input>
<ID>IN_1</ID>2525 </input>
<output>
<ID>OUT</ID>2520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2305</ID>
<type>AA_AND2</type>
<position>-1166,-3265</position>
<input>
<ID>IN_0</ID>2520 </input>
<input>
<ID>IN_1</ID>2527 </input>
<output>
<ID>OUT</ID>2521 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2306</ID>
<type>AA_AND2</type>
<position>-1294.5,-3192</position>
<input>
<ID>IN_0</ID>2503 </input>
<input>
<ID>IN_1</ID>2511 </input>
<output>
<ID>OUT</ID>2504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>2307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-759,-4532.5,-759,-4531.5</points>
<intersection>-4532.5 2</intersection>
<intersection>-4531.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-759,-4531.5,-581.5,-4531.5</points>
<connection>
<GID>1878</GID>
<name>N_in0</name></connection>
<intersection>-759 0</intersection>
<intersection>-581.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-764,-4532.5,-759,-4532.5</points>
<connection>
<GID>2031</GID>
<name>OUT</name></connection>
<intersection>-759 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-581.5,-4531.5,-581.5,-3636.5</points>
<connection>
<GID>2051</GID>
<name>IN_0</name></connection>
<intersection>-4531.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-785,-4550.5,-785,-4548</points>
<intersection>-4550.5 2</intersection>
<intersection>-4548 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-789,-4548,-785,-4548</points>
<connection>
<GID>2033</GID>
<name>Q</name></connection>
<intersection>-785 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-785,-4550.5,-781,-4550.5</points>
<connection>
<GID>2034</GID>
<name>IN_0</name></connection>
<intersection>-785 0</intersection></hsegment></shape></wire>
<wire>
<ID>2309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-845.5,-4713.5,-845.5,-4707.5</points>
<connection>
<GID>2417</GID>
<name>IN_0</name></connection>
<intersection>-4707.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-845.5,-4707.5,-777,-4707.5</points>
<connection>
<GID>2036</GID>
<name>OUT</name></connection>
<intersection>-845.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-770,-4706.5,-770,-4551.5</points>
<intersection>-4706.5 2</intersection>
<intersection>-4643.5 3</intersection>
<intersection>-4551.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-775,-4551.5,-770,-4551.5</points>
<connection>
<GID>2034</GID>
<name>OUT</name></connection>
<intersection>-770 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-771,-4706.5,-770,-4706.5</points>
<connection>
<GID>2036</GID>
<name>IN_1</name></connection>
<intersection>-770 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-770,-4643.5,-749.5,-4643.5</points>
<intersection>-770 0</intersection>
<intersection>-749.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-749.5,-4697,-749.5,-4643.5</points>
<intersection>-4697 5</intersection>
<intersection>-4687.5 11</intersection>
<intersection>-4679 13</intersection>
<intersection>-4670.5 15</intersection>
<intersection>-4663 17</intersection>
<intersection>-4643.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-760,-4697,-749.5,-4697</points>
<connection>
<GID>2038</GID>
<name>IN_1</name></connection>
<intersection>-749.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-760.5,-4687.5,-749.5,-4687.5</points>
<connection>
<GID>2040</GID>
<name>IN_1</name></connection>
<intersection>-749.5 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-760,-4679,-749.5,-4679</points>
<connection>
<GID>2042</GID>
<name>IN_1</name></connection>
<intersection>-749.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-760,-4670.5,-749.5,-4670.5</points>
<connection>
<GID>2044</GID>
<name>IN_1</name></connection>
<intersection>-749.5 4</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-759.5,-4663,-749.5,-4663</points>
<connection>
<GID>2046</GID>
<name>IN_1</name></connection>
<intersection>-749.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-832,-4713.5,-832,-4698</points>
<connection>
<GID>2418</GID>
<name>IN_0</name></connection>
<intersection>-4698 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-832,-4698,-766,-4698</points>
<connection>
<GID>2038</GID>
<name>OUT</name></connection>
<intersection>-832 0</intersection></hsegment></shape></wire>
<wire>
<ID>2312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-806,-4713.5,-806,-4680</points>
<connection>
<GID>2420</GID>
<name>IN_0</name></connection>
<intersection>-4680 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-806,-4680,-766,-4680</points>
<connection>
<GID>2042</GID>
<name>OUT</name></connection>
<intersection>-806 0</intersection></hsegment></shape></wire>
<wire>
<ID>2313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-793.5,-4714,-793.5,-4671.5</points>
<connection>
<GID>2421</GID>
<name>IN_0</name></connection>
<intersection>-4671.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-793.5,-4671.5,-766,-4671.5</points>
<connection>
<GID>2044</GID>
<name>OUT</name></connection>
<intersection>-793.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-781,-4714,-781,-4664</points>
<connection>
<GID>2423</GID>
<name>IN_0</name></connection>
<intersection>-4664 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-781,-4664,-765.5,-4664</points>
<connection>
<GID>2046</GID>
<name>OUT</name></connection>
<intersection>-781 0</intersection></hsegment></shape></wire>
<wire>
<ID>2315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-772,-4765.5,-772,-4764.5</points>
<intersection>-4765.5 1</intersection>
<intersection>-4764.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-775,-4765.5,-772,-4765.5</points>
<connection>
<GID>1883</GID>
<name>OUT</name></connection>
<intersection>-772 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-772,-4764.5,-768.5,-4764.5</points>
<connection>
<GID>2053</GID>
<name>IN_0</name></connection>
<intersection>-772 0</intersection></hsegment></shape></wire>
<wire>
<ID>2316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-803.5,-4782.5,-803.5,-4774.5</points>
<connection>
<GID>2416</GID>
<name>OUT</name></connection>
<intersection>-4782.5 8</intersection>
<intersection>-4776 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-803.5,-4776,-566.5,-4776</points>
<intersection>-803.5 0</intersection>
<intersection>-769 5</intersection>
<intersection>-566.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-566.5,-4776,-566.5,-3636.5</points>
<connection>
<GID>2055</GID>
<name>IN_1</name></connection>
<intersection>-4776 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-769,-4776,-769,-4766.5</points>
<intersection>-4776 1</intersection>
<intersection>-4766.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-769,-4766.5,-768.5,-4766.5</points>
<connection>
<GID>2053</GID>
<name>IN_1</name></connection>
<intersection>-769 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-803.5,-4782.5,-790.5,-4782.5</points>
<connection>
<GID>2056</GID>
<name>J</name></connection>
<intersection>-803.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-759.5,-4765.5,-759.5,-4765</points>
<intersection>-4765.5 2</intersection>
<intersection>-4765 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-759.5,-4765,-568.5,-4765</points>
<connection>
<GID>1886</GID>
<name>N_in0</name></connection>
<intersection>-759.5 0</intersection>
<intersection>-568.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-762.5,-4765.5,-759.5,-4765.5</points>
<connection>
<GID>2053</GID>
<name>OUT</name></connection>
<intersection>-759.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-568.5,-4765,-568.5,-3636.5</points>
<connection>
<GID>2055</GID>
<name>IN_0</name></connection>
<intersection>-4765 1</intersection></vsegment></shape></wire>
<wire>
<ID>2318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-780,-4788,-780,-4782.5</points>
<intersection>-4788 2</intersection>
<intersection>-4782.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-784.5,-4782.5,-780,-4782.5</points>
<connection>
<GID>2056</GID>
<name>Q</name></connection>
<intersection>-780 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-780,-4788,-775,-4788</points>
<connection>
<GID>2057</GID>
<name>IN_0</name></connection>
<intersection>-780 0</intersection></hsegment></shape></wire>
<wire>
<ID>2319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-836.5,-4940.5,-836.5,-4929</points>
<connection>
<GID>2456</GID>
<name>IN_0</name></connection>
<intersection>-4929 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-836.5,-4929,-759.5,-4929</points>
<connection>
<GID>2059</GID>
<name>OUT</name></connection>
<intersection>-836.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-750.5,-4928,-750.5,-4789</points>
<intersection>-4928 2</intersection>
<intersection>-4839.5 3</intersection>
<intersection>-4789 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-769,-4789,-750.5,-4789</points>
<connection>
<GID>2057</GID>
<name>OUT</name></connection>
<intersection>-750.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-753.5,-4928,-750.5,-4928</points>
<connection>
<GID>2059</GID>
<name>IN_1</name></connection>
<intersection>-750.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-750.5,-4839.5,-722.5,-4839.5</points>
<intersection>-750.5 0</intersection>
<intersection>-722.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-722.5,-4919.5,-722.5,-4839.5</points>
<intersection>-4919.5 5</intersection>
<intersection>-4909.5 7</intersection>
<intersection>-4900 9</intersection>
<intersection>-4891.5 11</intersection>
<intersection>-4883 13</intersection>
<intersection>-4839.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-741.5,-4919.5,-722.5,-4919.5</points>
<connection>
<GID>2062</GID>
<name>IN_1</name></connection>
<intersection>-722.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-740,-4909.5,-722.5,-4909.5</points>
<connection>
<GID>2064</GID>
<name>IN_1</name></connection>
<intersection>-722.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-739.5,-4900,-722.5,-4900</points>
<connection>
<GID>2118</GID>
<name>IN_1</name></connection>
<intersection>-722.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-740,-4891.5,-722.5,-4891.5</points>
<connection>
<GID>2125</GID>
<name>IN_1</name></connection>
<intersection>-722.5 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-740.5,-4883,-722.5,-4883</points>
<connection>
<GID>2303</GID>
<name>IN_1</name></connection>
<intersection>-722.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-823,-4940.5,-823,-4920.5</points>
<connection>
<GID>2457</GID>
<name>IN_0</name></connection>
<intersection>-4920.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-823,-4920.5,-747.5,-4920.5</points>
<connection>
<GID>2062</GID>
<name>OUT</name></connection>
<intersection>-823 0</intersection></hsegment></shape></wire>
<wire>
<ID>2322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-810,-4940.5,-810,-4910.5</points>
<connection>
<GID>2458</GID>
<name>IN_0</name></connection>
<intersection>-4910.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-810,-4910.5,-746,-4910.5</points>
<connection>
<GID>2064</GID>
<name>OUT</name></connection>
<intersection>-810 0</intersection></hsegment></shape></wire>
<wire>
<ID>2323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-797,-4940.5,-797,-4901</points>
<connection>
<GID>2459</GID>
<name>IN_0</name></connection>
<intersection>-4901 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-797,-4901,-745.5,-4901</points>
<connection>
<GID>2118</GID>
<name>OUT</name></connection>
<intersection>-797 0</intersection></hsegment></shape></wire>
<wire>
<ID>2324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-784.5,-4941,-784.5,-4892.5</points>
<connection>
<GID>2460</GID>
<name>IN_0</name></connection>
<intersection>-4892.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-784.5,-4892.5,-746,-4892.5</points>
<connection>
<GID>2125</GID>
<name>OUT</name></connection>
<intersection>-784.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-772,-4941,-772,-4884</points>
<connection>
<GID>2461</GID>
<name>IN_0</name></connection>
<intersection>-4884 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-772,-4884,-746.5,-4884</points>
<connection>
<GID>2303</GID>
<name>OUT</name></connection>
<intersection>-772 0</intersection></hsegment></shape></wire>
<wire>
<ID>2326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-763.5,-4992.5,-763.5,-4992</points>
<intersection>-4992.5 1</intersection>
<intersection>-4992 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-766,-4992.5,-763.5,-4992.5</points>
<connection>
<GID>1893</GID>
<name>OUT</name></connection>
<intersection>-763.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-763.5,-4992,-760.5,-4992</points>
<connection>
<GID>2361</GID>
<name>IN_0</name></connection>
<intersection>-763.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-935.5,-4022.5,-876.5,-4022.5</points>
<connection>
<GID>2025</GID>
<name>OUT</name></connection>
<connection>
<GID>2017</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-794.5,-5001.5,-553,-5001.5</points>
<connection>
<GID>2455</GID>
<name>OUT</name></connection>
<intersection>-762.5 5</intersection>
<intersection>-553 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-553,-5001.5,-553,-3175.5</points>
<intersection>-5001.5 1</intersection>
<intersection>-3637 9</intersection>
<intersection>-3175.5 7</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-762.5,-5001.5,-762.5,-4994</points>
<intersection>-5001.5 1</intersection>
<intersection>-4994 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-762.5,-4994,-760.5,-4994</points>
<connection>
<GID>2361</GID>
<name>IN_1</name></connection>
<intersection>-762.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1357.5,-3175.5,-553,-3175.5</points>
<intersection>-1357.5 8</intersection>
<intersection>-553 2</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-1357.5,-3190,-1357.5,-3175.5</points>
<connection>
<GID>2032</GID>
<name>IN_0</name></connection>
<intersection>-3175.5 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-554.5,-3637,-553,-3637</points>
<connection>
<GID>2422</GID>
<name>IN_1</name></connection>
<intersection>-553 2</intersection></hsegment></shape></wire>
<wire>
<ID>2329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-754.5,-4993,-556.5,-4993</points>
<connection>
<GID>2361</GID>
<name>OUT</name></connection>
<connection>
<GID>1891</GID>
<name>N_in0</name></connection>
<intersection>-556.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-556.5,-4993,-556.5,-3637</points>
<connection>
<GID>2422</GID>
<name>IN_0</name></connection>
<intersection>-4993 1</intersection></vsegment></shape></wire>
<wire>
<ID>2330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-594.5,-3630.5,-594.5,-3624</points>
<connection>
<GID>1987</GID>
<name>OUT</name></connection>
<intersection>-3624 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-578.5,-3624,-578.5,-3618</points>
<connection>
<GID>2425</GID>
<name>IN_0</name></connection>
<intersection>-3624 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-594.5,-3624,-578.5,-3624</points>
<intersection>-594.5 0</intersection>
<intersection>-578.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-580.5,-3630.5,-580.5,-3625</points>
<connection>
<GID>2051</GID>
<name>OUT</name></connection>
<intersection>-3625 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-576.5,-3625,-576.5,-3618</points>
<connection>
<GID>2425</GID>
<name>IN_1</name></connection>
<intersection>-3625 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-580.5,-3625,-576.5,-3625</points>
<intersection>-580.5 0</intersection>
<intersection>-576.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-567.5,-3630.5,-567.5,-3624</points>
<connection>
<GID>2055</GID>
<name>OUT</name></connection>
<intersection>-3624 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-574.5,-3624,-574.5,-3618</points>
<connection>
<GID>2425</GID>
<name>IN_2</name></connection>
<intersection>-3624 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-574.5,-3624,-567.5,-3624</points>
<intersection>-574.5 1</intersection>
<intersection>-567.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-555.5,-3631,-555.5,-3622</points>
<connection>
<GID>2422</GID>
<name>OUT</name></connection>
<intersection>-3622 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-572.5,-3622,-572.5,-3618</points>
<connection>
<GID>2425</GID>
<name>IN_3</name></connection>
<intersection>-3622 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-572.5,-3622,-555.5,-3622</points>
<intersection>-572.5 1</intersection>
<intersection>-555.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-640.5,-3613.5,-640.5,-3604.5</points>
<connection>
<GID>1866</GID>
<name>OUT</name></connection>
<intersection>-3604.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-614.5,-3604.5,-614.5,-3596</points>
<connection>
<GID>2462</GID>
<name>IN_0</name></connection>
<intersection>-3604.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-640.5,-3604.5,-614.5,-3604.5</points>
<intersection>-640.5 0</intersection>
<intersection>-614.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-612.5,-3604,-612.5,-3596</points>
<connection>
<GID>2462</GID>
<name>IN_1</name></connection>
<intersection>-3604 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-575.5,-3612,-575.5,-3604</points>
<connection>
<GID>2425</GID>
<name>OUT</name></connection>
<intersection>-3604 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-612.5,-3604,-575.5,-3604</points>
<intersection>-612.5 0</intersection>
<intersection>-575.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-853.5,-4058.5,-853.5,-4022.5</points>
<connection>
<GID>2008</GID>
<name>IN_1</name></connection>
<intersection>-4022.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-870.5,-4022.5,-853.5,-4022.5</points>
<connection>
<GID>2017</GID>
<name>Q</name></connection>
<intersection>-853.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2337</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-936,-4012.5,-889.5,-4012.5</points>
<connection>
<GID>2026</GID>
<name>OUT</name></connection>
<connection>
<GID>2018</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-840,-4058.5,-840,-4012.5</points>
<connection>
<GID>2009</GID>
<name>IN_1</name></connection>
<intersection>-4012.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-883.5,-4012.5,-840,-4012.5</points>
<connection>
<GID>2018</GID>
<name>Q</name></connection>
<intersection>-840 0</intersection></hsegment></shape></wire>
<wire>
<ID>2339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-937.5,-4001.5,-902.5,-4001.5</points>
<connection>
<GID>2027</GID>
<name>OUT</name></connection>
<connection>
<GID>2019</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-827,-4058.5,-827,-4001.5</points>
<connection>
<GID>2010</GID>
<name>IN_1</name></connection>
<intersection>-4001.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-896.5,-4001.5,-827,-4001.5</points>
<connection>
<GID>2019</GID>
<name>Q</name></connection>
<intersection>-827 0</intersection></hsegment></shape></wire>
<wire>
<ID>2341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-938,-3992.5,-910,-3992.5</points>
<connection>
<GID>2028</GID>
<name>OUT</name></connection>
<connection>
<GID>2021</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-814,-4058.5,-814,-3992.5</points>
<connection>
<GID>2011</GID>
<name>IN_1</name></connection>
<intersection>-3992.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-904,-3992.5,-814,-3992.5</points>
<connection>
<GID>2021</GID>
<name>Q</name></connection>
<intersection>-814 0</intersection></hsegment></shape></wire>
<wire>
<ID>2343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-939,-3985,-918.5,-3985</points>
<connection>
<GID>2039</GID>
<name>OUT</name></connection>
<connection>
<GID>2022</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-801.5,-4059,-801.5,-3985</points>
<connection>
<GID>2012</GID>
<name>IN_1</name></connection>
<intersection>-3985 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-912.5,-3985,-801.5,-3985</points>
<connection>
<GID>2022</GID>
<name>Q</name></connection>
<intersection>-801.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-940,-3977.5,-927.5,-3977.5</points>
<connection>
<GID>2067</GID>
<name>OUT</name></connection>
<connection>
<GID>2023</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-789,-4059,-789,-3977.5</points>
<connection>
<GID>2014</GID>
<name>IN_1</name></connection>
<intersection>-3977.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-921.5,-3977.5,-789,-3977.5</points>
<connection>
<GID>2023</GID>
<name>Q</name></connection>
<intersection>-789 0</intersection></hsegment></shape></wire>
<wire>
<ID>2347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-933,-4024.5,-933,-3973.5</points>
<connection>
<GID>2024</GID>
<name>OUT_0</name></connection>
<intersection>-4024.5 7</intersection>
<intersection>-4014.5 5</intersection>
<intersection>-4003.5 8</intersection>
<intersection>-3994.5 3</intersection>
<intersection>-3987 9</intersection>
<intersection>-3979.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-933,-3979.5,-927.5,-3979.5</points>
<connection>
<GID>2023</GID>
<name>clock</name></connection>
<intersection>-933 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-933,-3994.5,-910,-3994.5</points>
<connection>
<GID>2021</GID>
<name>clock</name></connection>
<intersection>-933 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-933,-4014.5,-889.5,-4014.5</points>
<connection>
<GID>2018</GID>
<name>clock</name></connection>
<intersection>-933 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-933,-4024.5,-876.5,-4024.5</points>
<connection>
<GID>2017</GID>
<name>clock</name></connection>
<intersection>-933 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-933,-4003.5,-902.5,-4003.5</points>
<connection>
<GID>2019</GID>
<name>clock</name></connection>
<intersection>-933 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-933,-3987,-918.5,-3987</points>
<connection>
<GID>2022</GID>
<name>clock</name></connection>
<intersection>-933 0</intersection></hsegment></shape></wire>
<wire>
<ID>2348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-611.5,-3431,-611.5,-3272.5</points>
<intersection>-3431 2</intersection>
<intersection>-3272.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-613.5,-3590,-613.5,-3431</points>
<connection>
<GID>2462</GID>
<name>OUT</name></connection>
<intersection>-3431 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-613.5,-3431,-611.5,-3431</points>
<intersection>-613.5 1</intersection>
<intersection>-611.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1091.5,-3272.5,-611.5,-3272.5</points>
<connection>
<GID>2257</GID>
<name>clear</name></connection>
<intersection>-611.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-961.5,-4310.5,-961.5,-4157</points>
<intersection>-4310.5 13</intersection>
<intersection>-4220.5 1</intersection>
<intersection>-4210.5 3</intersection>
<intersection>-4199.5 5</intersection>
<intersection>-4190.5 7</intersection>
<intersection>-4183 9</intersection>
<intersection>-4157 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-961.5,-4220.5,-931,-4220.5</points>
<connection>
<GID>2141</GID>
<name>IN_0</name></connection>
<intersection>-961.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-961.5,-4210.5,-931.5,-4210.5</points>
<connection>
<GID>2143</GID>
<name>IN_0</name></connection>
<intersection>-961.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-961.5,-4199.5,-933,-4199.5</points>
<connection>
<GID>2145</GID>
<name>IN_0</name></connection>
<intersection>-961.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-961.5,-4190.5,-933.5,-4190.5</points>
<connection>
<GID>2147</GID>
<name>IN_0</name></connection>
<intersection>-961.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-961.5,-4183,-934.5,-4183</points>
<connection>
<GID>2149</GID>
<name>IN_0</name></connection>
<intersection>-961.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-961.5,-4157,-797.5,-4157</points>
<intersection>-961.5 0</intersection>
<intersection>-961 17</intersection>
<intersection>-935.5 16</intersection>
<intersection>-797.5 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-961.5,-4310.5,-778,-4310.5</points>
<connection>
<GID>1876</GID>
<name>IN_1</name></connection>
<intersection>-961.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-797.5,-4157,-797.5,-4139</points>
<intersection>-4157 11</intersection>
<intersection>-4139 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-797.5,-4139,-788,-4139</points>
<connection>
<GID>1969</GID>
<name>IN_1</name></connection>
<intersection>-797.5 14</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-935.5,-4175.5,-935.5,-4157</points>
<connection>
<GID>2151</GID>
<name>IN_0</name></connection>
<intersection>-4157 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-961,-4157,-961,-4152</points>
<connection>
<GID>2105</GID>
<name>OUT</name></connection>
<intersection>-4157 11</intersection></vsegment></shape></wire>
<wire>
<ID>2350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-842,-4267,-842,-4263.5</points>
<connection>
<GID>2107</GID>
<name>OUT</name></connection>
<intersection>-4267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-842,-4267,-841,-4267</points>
<connection>
<GID>2153</GID>
<name>IN_0</name></connection>
<intersection>-842 0</intersection></hsegment></shape></wire>
<wire>
<ID>2351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-828.5,-4267.5,-828.5,-4263.5</points>
<connection>
<GID>2110</GID>
<name>OUT</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-828.5,-4267.5,-825,-4267.5</points>
<connection>
<GID>2070</GID>
<name>IN_0</name></connection>
<intersection>-828.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-815.5,-4267.5,-815.5,-4263.5</points>
<connection>
<GID>2112</GID>
<name>OUT</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-815.5,-4267.5,-811.5,-4267.5</points>
<connection>
<GID>2072</GID>
<name>IN_0</name></connection>
<intersection>-815.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-799.5,-4267.5,-799.5,-4263.5</points>
<intersection>-4267.5 1</intersection>
<intersection>-4263.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-799.5,-4267.5,-796.5,-4267.5</points>
<connection>
<GID>2073</GID>
<name>IN_0</name></connection>
<intersection>-799.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-802.5,-4263.5,-799.5,-4263.5</points>
<connection>
<GID>2114</GID>
<name>OUT</name></connection>
<intersection>-799.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-790,-4266,-790,-4264</points>
<connection>
<GID>2116</GID>
<name>OUT</name></connection>
<intersection>-4266 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-790,-4266,-786,-4266</points>
<intersection>-790 0</intersection>
<intersection>-786 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-786,-4267.5,-786,-4266</points>
<connection>
<GID>2075</GID>
<name>IN_0</name></connection>
<intersection>-4266 1</intersection></vsegment></shape></wire>
<wire>
<ID>2355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-777.5,-4266,-777.5,-4264</points>
<connection>
<GID>2120</GID>
<name>OUT</name></connection>
<intersection>-4266 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-777.5,-4266,-773,-4266</points>
<intersection>-777.5 0</intersection>
<intersection>-773 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-773,-4267.5,-773,-4266</points>
<connection>
<GID>2076</GID>
<name>IN_0</name></connection>
<intersection>-4266 1</intersection></vsegment></shape></wire>
<wire>
<ID>2356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-831,-4275,-831,-4267</points>
<connection>
<GID>2078</GID>
<name>IN_0</name></connection>
<intersection>-4267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-835,-4267,-831,-4267</points>
<connection>
<GID>2153</GID>
<name>OUT_0</name></connection>
<intersection>-831 0</intersection></hsegment></shape></wire>
<wire>
<ID>2357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-816,-4275,-816,-4267.5</points>
<connection>
<GID>2079</GID>
<name>IN_0</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-819,-4267.5,-816,-4267.5</points>
<connection>
<GID>2070</GID>
<name>OUT_0</name></connection>
<intersection>-816 0</intersection></hsegment></shape></wire>
<wire>
<ID>2358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-801,-4275,-801,-4267.5</points>
<connection>
<GID>2081</GID>
<name>IN_0</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-805.5,-4267.5,-801,-4267.5</points>
<connection>
<GID>2072</GID>
<name>OUT_0</name></connection>
<intersection>-801 0</intersection></hsegment></shape></wire>
<wire>
<ID>2359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-789.5,-4274.5,-789.5,-4267.5</points>
<connection>
<GID>2083</GID>
<name>IN_0</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-790.5,-4267.5,-789.5,-4267.5</points>
<connection>
<GID>2073</GID>
<name>OUT_0</name></connection>
<intersection>-789.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776.5,-4275,-776.5,-4267.5</points>
<connection>
<GID>2085</GID>
<name>IN_0</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-780,-4267.5,-776.5,-4267.5</points>
<connection>
<GID>2075</GID>
<name>OUT_0</name></connection>
<intersection>-776.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-763.5,-4274.5,-763.5,-4267.5</points>
<connection>
<GID>2087</GID>
<name>IN_0</name></connection>
<intersection>-4267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-767,-4267.5,-763.5,-4267.5</points>
<connection>
<GID>2076</GID>
<name>OUT_0</name></connection>
<intersection>-763.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-831,-4284.5,-831,-4279</points>
<connection>
<GID>2078</GID>
<name>OUT_0</name></connection>
<intersection>-4284.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-816,-4290.5,-816,-4284.5</points>
<connection>
<GID>2091</GID>
<name>IN_3</name></connection>
<intersection>-4284.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-831,-4284.5,-816,-4284.5</points>
<intersection>-831 0</intersection>
<intersection>-816 1</intersection></hsegment></shape></wire>
<wire>
<ID>2363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-816,-4284,-816,-4279</points>
<connection>
<GID>2079</GID>
<name>OUT_0</name></connection>
<intersection>-4284 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-814,-4290.5,-814,-4284</points>
<connection>
<GID>2091</GID>
<name>IN_2</name></connection>
<intersection>-4284 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-816,-4284,-814,-4284</points>
<intersection>-816 0</intersection>
<intersection>-814 1</intersection></hsegment></shape></wire>
<wire>
<ID>2364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-801,-4284.5,-801,-4279</points>
<connection>
<GID>2081</GID>
<name>OUT_0</name></connection>
<intersection>-4284.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-812,-4290.5,-812,-4284.5</points>
<connection>
<GID>2091</GID>
<name>IN_1</name></connection>
<intersection>-4284.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-812,-4284.5,-801,-4284.5</points>
<intersection>-812 1</intersection>
<intersection>-801 0</intersection></hsegment></shape></wire>
<wire>
<ID>2365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-789.5,-4285.5,-789.5,-4278.5</points>
<connection>
<GID>2083</GID>
<name>OUT_0</name></connection>
<intersection>-4285.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-810,-4290.5,-810,-4285.5</points>
<connection>
<GID>2091</GID>
<name>IN_0</name></connection>
<intersection>-4285.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-810,-4285.5,-789.5,-4285.5</points>
<intersection>-810 1</intersection>
<intersection>-789.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776.5,-4284,-776.5,-4279</points>
<connection>
<GID>2085</GID>
<name>OUT_0</name></connection>
<intersection>-4284 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-777.5,-4289.5,-777.5,-4284</points>
<connection>
<GID>2099</GID>
<name>IN_1</name></connection>
<intersection>-4284 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-777.5,-4284,-776.5,-4284</points>
<intersection>-777.5 1</intersection>
<intersection>-776.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-763.5,-4284,-763.5,-4278.5</points>
<connection>
<GID>2087</GID>
<name>OUT_0</name></connection>
<intersection>-4284 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-775.5,-4289.5,-775.5,-4284</points>
<connection>
<GID>2099</GID>
<name>IN_0</name></connection>
<intersection>-4284 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-775.5,-4284,-763.5,-4284</points>
<intersection>-775.5 1</intersection>
<intersection>-763.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-813,-4299.5,-813,-4296.5</points>
<connection>
<GID>2091</GID>
<name>OUT</name></connection>
<intersection>-4299.5 2</intersection>
<intersection>-4299 8</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-800,-4312.5,-800,-4299.5</points>
<connection>
<GID>2103</GID>
<name>IN_1</name></connection>
<intersection>-4307.5 7</intersection>
<intersection>-4299.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-813,-4299.5,-800,-4299.5</points>
<intersection>-813 0</intersection>
<intersection>-800 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-800,-4307.5,-788.5,-4307.5</points>
<connection>
<GID>2133</GID>
<name>IN_0</name></connection>
<intersection>-800 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-868.5,-4299,-813,-4299</points>
<connection>
<GID>1901</GID>
<name>IN_0</name></connection>
<intersection>-813 0</intersection></hsegment></shape></wire>
<wire>
<ID>2369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776.5,-4299,-776.5,-4295.5</points>
<connection>
<GID>2099</GID>
<name>OUT</name></connection>
<intersection>-4299 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-798,-4312.5,-798,-4299</points>
<connection>
<GID>2103</GID>
<name>IN_0</name></connection>
<intersection>-4309.5 6</intersection>
<intersection>-4303.5 7</intersection>
<intersection>-4299 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-798,-4299,-776.5,-4299</points>
<intersection>-798 1</intersection>
<intersection>-776.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-798,-4309.5,-788.5,-4309.5</points>
<connection>
<GID>2133</GID>
<name>IN_1</name></connection>
<intersection>-798 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-909,-4303.5,-798,-4303.5</points>
<intersection>-909 8</intersection>
<intersection>-798 1</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-909,-4303.5,-909,-4301</points>
<connection>
<GID>1895</GID>
<name>IN_0</name></connection>
<intersection>-4303.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>2370</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-925,-4221.5,-866,-4221.5</points>
<connection>
<GID>2141</GID>
<name>OUT</name></connection>
<connection>
<GID>2127</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-843,-4257.5,-843,-4221.5</points>
<connection>
<GID>2107</GID>
<name>IN_1</name></connection>
<intersection>-4221.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-860,-4221.5,-843,-4221.5</points>
<connection>
<GID>2127</GID>
<name>Q</name></connection>
<intersection>-843 0</intersection></hsegment></shape></wire>
<wire>
<ID>2372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-925.5,-4211.5,-879,-4211.5</points>
<connection>
<GID>2143</GID>
<name>OUT</name></connection>
<connection>
<GID>2129</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-829.5,-4257.5,-829.5,-4211.5</points>
<connection>
<GID>2110</GID>
<name>IN_1</name></connection>
<intersection>-4211.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-873,-4211.5,-829.5,-4211.5</points>
<connection>
<GID>2129</GID>
<name>Q</name></connection>
<intersection>-829.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-927,-4200.5,-892,-4200.5</points>
<connection>
<GID>2145</GID>
<name>OUT</name></connection>
<connection>
<GID>2131</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-816.5,-4257.5,-816.5,-4200.5</points>
<connection>
<GID>2112</GID>
<name>IN_1</name></connection>
<intersection>-4200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-886,-4200.5,-816.5,-4200.5</points>
<connection>
<GID>2131</GID>
<name>Q</name></connection>
<intersection>-816.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-927.5,-4191.5,-899.5,-4191.5</points>
<connection>
<GID>2147</GID>
<name>OUT</name></connection>
<connection>
<GID>2135</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-803.5,-4257.5,-803.5,-4191.5</points>
<connection>
<GID>2114</GID>
<name>IN_1</name></connection>
<intersection>-4191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-893.5,-4191.5,-803.5,-4191.5</points>
<connection>
<GID>2135</GID>
<name>Q</name></connection>
<intersection>-803.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2378</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-928.5,-4184,-908,-4184</points>
<connection>
<GID>2149</GID>
<name>OUT</name></connection>
<connection>
<GID>2137</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-791,-4258,-791,-4184</points>
<connection>
<GID>2116</GID>
<name>IN_1</name></connection>
<intersection>-4184 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-902,-4184,-791,-4184</points>
<connection>
<GID>2137</GID>
<name>Q</name></connection>
<intersection>-791 0</intersection></hsegment></shape></wire>
<wire>
<ID>2380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-929.5,-4176.5,-917,-4176.5</points>
<connection>
<GID>2151</GID>
<name>OUT</name></connection>
<connection>
<GID>2138</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-778.5,-4258,-778.5,-4176.5</points>
<connection>
<GID>2120</GID>
<name>IN_1</name></connection>
<intersection>-4176.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-911,-4176.5,-778.5,-4176.5</points>
<connection>
<GID>2138</GID>
<name>Q</name></connection>
<intersection>-778.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-922,-4223.5,-922,-4172.5</points>
<connection>
<GID>2140</GID>
<name>OUT_0</name></connection>
<intersection>-4223.5 7</intersection>
<intersection>-4213.5 5</intersection>
<intersection>-4202.5 8</intersection>
<intersection>-4193.5 3</intersection>
<intersection>-4186 9</intersection>
<intersection>-4178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-922,-4178.5,-917,-4178.5</points>
<connection>
<GID>2138</GID>
<name>clock</name></connection>
<intersection>-922 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-922,-4193.5,-899.5,-4193.5</points>
<connection>
<GID>2135</GID>
<name>clock</name></connection>
<intersection>-922 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-922,-4213.5,-879,-4213.5</points>
<connection>
<GID>2129</GID>
<name>clock</name></connection>
<intersection>-922 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-922,-4223.5,-866,-4223.5</points>
<connection>
<GID>2127</GID>
<name>clock</name></connection>
<intersection>-922 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-922,-4202.5,-892,-4202.5</points>
<connection>
<GID>2131</GID>
<name>clock</name></connection>
<intersection>-922 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-922,-4186,-908,-4186</points>
<connection>
<GID>2137</GID>
<name>clock</name></connection>
<intersection>-922 0</intersection></hsegment></shape></wire>
<wire>
<ID>2383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805,-3741,-805,-3736</points>
<connection>
<GID>1928</GID>
<name>OUT_0</name></connection>
<intersection>-3741 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-806,-3746.5,-806,-3741</points>
<connection>
<GID>2160</GID>
<name>IN_1</name></connection>
<intersection>-3741 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-806,-3741,-805,-3741</points>
<intersection>-806 1</intersection>
<intersection>-805 0</intersection></hsegment></shape></wire>
<wire>
<ID>2384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-792,-3741,-792,-3735.5</points>
<connection>
<GID>1929</GID>
<name>OUT_0</name></connection>
<intersection>-3741 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-804,-3746.5,-804,-3741</points>
<connection>
<GID>2160</GID>
<name>IN_0</name></connection>
<intersection>-3741 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-804,-3741,-792,-3741</points>
<intersection>-804 1</intersection>
<intersection>-792 0</intersection></hsegment></shape></wire>
<wire>
<ID>2385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-841.5,-3756.5,-841.5,-3753.5</points>
<connection>
<GID>2159</GID>
<name>OUT</name></connection>
<intersection>-3756.5 2</intersection>
<intersection>-3753.5 5</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-827,-3764.5,-827,-3756.5</points>
<connection>
<GID>2161</GID>
<name>IN_1</name></connection>
<intersection>-3758.5 3</intersection>
<intersection>-3756.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-841.5,-3756.5,-827,-3756.5</points>
<intersection>-841.5 0</intersection>
<intersection>-827 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-827,-3758.5,-788.5,-3758.5</points>
<connection>
<GID>1865</GID>
<name>IN_1</name></connection>
<intersection>-827 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-861.5,-3753.5,-841.5,-3753.5</points>
<intersection>-861.5 6</intersection>
<intersection>-841.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-861.5,-3754,-861.5,-3753.5</points>
<intersection>-3754 10</intersection>
<intersection>-3753.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-949.5,-3754,-861.5,-3754</points>
<connection>
<GID>2054</GID>
<name>IN_0</name></connection>
<intersection>-861.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>2386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805,-3756.5,-805,-3752.5</points>
<connection>
<GID>2160</GID>
<name>OUT</name></connection>
<intersection>-3756.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-825,-3764.5,-825,-3756.5</points>
<connection>
<GID>2161</GID>
<name>IN_0</name></connection>
<intersection>-3759.5 4</intersection>
<intersection>-3756.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-825,-3756.5,-788.5,-3756.5</points>
<connection>
<GID>1865</GID>
<name>IN_0</name></connection>
<intersection>-825 1</intersection>
<intersection>-805 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-959.5,-3759.5,-825,-3759.5</points>
<intersection>-959.5 5</intersection>
<intersection>-825 1</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-959.5,-3759.5,-959.5,-3755</points>
<intersection>-3759.5 4</intersection>
<intersection>-3755 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-961.5,-3755,-959.5,-3755</points>
<connection>
<GID>2049</GID>
<name>IN_0</name></connection>
<intersection>-959.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>2387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-967.5,-4532.5,-967.5,-4369.5</points>
<connection>
<GID>2115</GID>
<name>OUT</name></connection>
<intersection>-4532.5 13</intersection>
<intersection>-4442.5 1</intersection>
<intersection>-4432.5 3</intersection>
<intersection>-4421.5 5</intersection>
<intersection>-4412.5 7</intersection>
<intersection>-4405 9</intersection>
<intersection>-4373 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-967.5,-4442.5,-937.5,-4442.5</points>
<connection>
<GID>2394</GID>
<name>IN_0</name></connection>
<intersection>-967.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-967.5,-4432.5,-938,-4432.5</points>
<connection>
<GID>2396</GID>
<name>IN_0</name></connection>
<intersection>-967.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-967.5,-4421.5,-939.5,-4421.5</points>
<connection>
<GID>2397</GID>
<name>IN_0</name></connection>
<intersection>-967.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-967.5,-4412.5,-940,-4412.5</points>
<connection>
<GID>2398</GID>
<name>IN_0</name></connection>
<intersection>-967.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-967.5,-4405,-941,-4405</points>
<connection>
<GID>2399</GID>
<name>IN_0</name></connection>
<intersection>-967.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-967.5,-4373,-775,-4373</points>
<intersection>-967.5 0</intersection>
<intersection>-942 15</intersection>
<intersection>-775 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-967.5,-4532.5,-782.5,-4532.5</points>
<connection>
<GID>1880</GID>
<name>IN_1</name></connection>
<intersection>-967.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-775,-4373,-775,-4334.5</points>
<connection>
<GID>1990</GID>
<name>IN_1</name></connection>
<intersection>-4373 11</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-942,-4397.5,-942,-4373</points>
<connection>
<GID>2400</GID>
<name>IN_0</name></connection>
<intersection>-4373 11</intersection></vsegment></shape></wire>
<wire>
<ID>2388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-848.5,-4489,-848.5,-4485.5</points>
<connection>
<GID>2352</GID>
<name>OUT</name></connection>
<intersection>-4489 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-848.5,-4489,-847.5,-4489</points>
<connection>
<GID>2401</GID>
<name>IN_0</name></connection>
<intersection>-848.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-835,-4489.5,-835,-4485.5</points>
<connection>
<GID>2354</GID>
<name>OUT</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-835,-4489.5,-831.5,-4489.5</points>
<connection>
<GID>2155</GID>
<name>IN_0</name></connection>
<intersection>-835 0</intersection></hsegment></shape></wire>
<wire>
<ID>2390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-822,-4489.5,-822,-4485.5</points>
<connection>
<GID>2356</GID>
<name>OUT</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-822,-4489.5,-817.5,-4489.5</points>
<connection>
<GID>2156</GID>
<name>IN_0</name></connection>
<intersection>-822 0</intersection></hsegment></shape></wire>
<wire>
<ID>2391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-806,-4489.5,-806,-4485.5</points>
<intersection>-4489.5 1</intersection>
<intersection>-4485.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-806,-4489.5,-803,-4489.5</points>
<connection>
<GID>2157</GID>
<name>IN_0</name></connection>
<intersection>-806 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-809,-4485.5,-806,-4485.5</points>
<connection>
<GID>2357</GID>
<name>OUT</name></connection>
<intersection>-806 0</intersection></hsegment></shape></wire>
<wire>
<ID>2392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-796.5,-4488,-796.5,-4486</points>
<connection>
<GID>2358</GID>
<name>OUT</name></connection>
<intersection>-4488 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-796.5,-4488,-792.5,-4488</points>
<intersection>-796.5 0</intersection>
<intersection>-792.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-792.5,-4489.5,-792.5,-4488</points>
<connection>
<GID>2158</GID>
<name>IN_0</name></connection>
<intersection>-4488 1</intersection></vsegment></shape></wire>
<wire>
<ID>2393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-990,-3552.5,-990,-3503</points>
<connection>
<GID>2071</GID>
<name>OUT</name></connection>
<intersection>-3552.5 1</intersection>
<intersection>-3542.5 3</intersection>
<intersection>-3531.5 5</intersection>
<intersection>-3522.5 7</intersection>
<intersection>-3515 9</intersection>
<intersection>-3507.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-990,-3552.5,-959,-3552.5</points>
<connection>
<GID>2171</GID>
<name>IN_0</name></connection>
<intersection>-990 0</intersection>
<intersection>-974.5 12</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-990,-3542.5,-959.5,-3542.5</points>
<connection>
<GID>2174</GID>
<name>IN_0</name></connection>
<intersection>-990 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-990,-3531.5,-961,-3531.5</points>
<connection>
<GID>2175</GID>
<name>IN_0</name></connection>
<intersection>-990 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-990,-3522.5,-961.5,-3522.5</points>
<connection>
<GID>2177</GID>
<name>IN_0</name></connection>
<intersection>-990 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-990,-3515,-962.5,-3515</points>
<connection>
<GID>2180</GID>
<name>IN_0</name></connection>
<intersection>-990 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-990,-3507.5,-963.5,-3507.5</points>
<connection>
<GID>2181</GID>
<name>IN_0</name></connection>
<intersection>-990 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-974.5,-3648.5,-974.5,-3552.5</points>
<intersection>-3648.5 13</intersection>
<intersection>-3552.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-974.5,-3648.5,-793.5,-3648.5</points>
<intersection>-974.5 12</intersection>
<intersection>-793.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-793.5,-3648.5,-793.5,-3648</points>
<connection>
<GID>1861</GID>
<name>IN_1</name></connection>
<intersection>-3648.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>2394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-784,-4488,-784,-4486</points>
<connection>
<GID>2359</GID>
<name>OUT</name></connection>
<intersection>-4488 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-784,-4488,-779.5,-4488</points>
<intersection>-784 0</intersection>
<intersection>-779.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-779.5,-4489.5,-779.5,-4488</points>
<connection>
<GID>2169</GID>
<name>IN_0</name></connection>
<intersection>-4488 1</intersection></vsegment></shape></wire>
<wire>
<ID>2395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-837.5,-4497,-837.5,-4489</points>
<connection>
<GID>2170</GID>
<name>IN_0</name></connection>
<intersection>-4489 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-841.5,-4489,-837.5,-4489</points>
<connection>
<GID>2401</GID>
<name>OUT_0</name></connection>
<intersection>-837.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-870,-3599,-870,-3595.5</points>
<connection>
<GID>2331</GID>
<name>OUT</name></connection>
<intersection>-3599 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-870,-3599,-869,-3599</points>
<connection>
<GID>2196</GID>
<name>IN_0</name></connection>
<intersection>-870 0</intersection></hsegment></shape></wire>
<wire>
<ID>2397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-856.5,-3599.5,-856.5,-3595.5</points>
<connection>
<GID>2332</GID>
<name>OUT</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-856.5,-3599.5,-853,-3599.5</points>
<connection>
<GID>2221</GID>
<name>IN_0</name></connection>
<intersection>-856.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-843.5,-3599.5,-843.5,-3595.5</points>
<connection>
<GID>2334</GID>
<name>OUT</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-843.5,-3599.5,-839.5,-3599.5</points>
<connection>
<GID>2230</GID>
<name>IN_0</name></connection>
<intersection>-843.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-827.5,-3599.5,-827.5,-3595.5</points>
<intersection>-3599.5 1</intersection>
<intersection>-3595.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-827.5,-3599.5,-824.5,-3599.5</points>
<connection>
<GID>2237</GID>
<name>IN_0</name></connection>
<intersection>-827.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-830.5,-3595.5,-827.5,-3595.5</points>
<connection>
<GID>2336</GID>
<name>OUT</name></connection>
<intersection>-827.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-818,-3598,-818,-3596</points>
<connection>
<GID>2337</GID>
<name>OUT</name></connection>
<intersection>-3598 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-818,-3598,-814,-3598</points>
<intersection>-818 0</intersection>
<intersection>-814 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-814,-3599.5,-814,-3598</points>
<connection>
<GID>2242</GID>
<name>IN_0</name></connection>
<intersection>-3598 1</intersection></vsegment></shape></wire>
<wire>
<ID>2401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805.5,-3598,-805.5,-3596</points>
<connection>
<GID>2339</GID>
<name>OUT</name></connection>
<intersection>-3598 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-805.5,-3598,-801,-3598</points>
<intersection>-805.5 0</intersection>
<intersection>-801 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-801,-3599.5,-801,-3598</points>
<connection>
<GID>2249</GID>
<name>IN_0</name></connection>
<intersection>-3598 1</intersection></vsegment></shape></wire>
<wire>
<ID>2402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-859,-3607,-859,-3599</points>
<connection>
<GID>2253</GID>
<name>IN_0</name></connection>
<intersection>-3599 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-863,-3599,-859,-3599</points>
<connection>
<GID>2196</GID>
<name>OUT_0</name></connection>
<intersection>-859 0</intersection></hsegment></shape></wire>
<wire>
<ID>2403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844,-3607,-844,-3599.5</points>
<connection>
<GID>2256</GID>
<name>IN_0</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-847,-3599.5,-844,-3599.5</points>
<connection>
<GID>2221</GID>
<name>OUT_0</name></connection>
<intersection>-844 0</intersection></hsegment></shape></wire>
<wire>
<ID>2404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-829,-3607,-829,-3599.5</points>
<connection>
<GID>2259</GID>
<name>IN_0</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-833.5,-3599.5,-829,-3599.5</points>
<connection>
<GID>2230</GID>
<name>OUT_0</name></connection>
<intersection>-829 0</intersection></hsegment></shape></wire>
<wire>
<ID>2405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-817.5,-3606.5,-817.5,-3599.5</points>
<connection>
<GID>2261</GID>
<name>IN_0</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-818.5,-3599.5,-817.5,-3599.5</points>
<connection>
<GID>2237</GID>
<name>OUT_0</name></connection>
<intersection>-817.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-804.5,-3607,-804.5,-3599.5</points>
<connection>
<GID>2263</GID>
<name>IN_0</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-808,-3599.5,-804.5,-3599.5</points>
<connection>
<GID>2242</GID>
<name>OUT_0</name></connection>
<intersection>-804.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-791.5,-3606.5,-791.5,-3599.5</points>
<connection>
<GID>2266</GID>
<name>IN_0</name></connection>
<intersection>-3599.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-795,-3599.5,-791.5,-3599.5</points>
<connection>
<GID>2249</GID>
<name>OUT_0</name></connection>
<intersection>-791.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-859,-3616.5,-859,-3611</points>
<connection>
<GID>2253</GID>
<name>OUT_0</name></connection>
<intersection>-3616.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-844,-3622.5,-844,-3616.5</points>
<connection>
<GID>2282</GID>
<name>IN_3</name></connection>
<intersection>-3616.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-859,-3616.5,-844,-3616.5</points>
<intersection>-859 0</intersection>
<intersection>-844 1</intersection></hsegment></shape></wire>
<wire>
<ID>2409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844,-3616,-844,-3611</points>
<connection>
<GID>2256</GID>
<name>OUT_0</name></connection>
<intersection>-3616 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-842,-3622.5,-842,-3616</points>
<connection>
<GID>2282</GID>
<name>IN_2</name></connection>
<intersection>-3616 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-844,-3616,-842,-3616</points>
<intersection>-844 0</intersection>
<intersection>-842 1</intersection></hsegment></shape></wire>
<wire>
<ID>2410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-829,-3616.5,-829,-3611</points>
<connection>
<GID>2259</GID>
<name>OUT_0</name></connection>
<intersection>-3616.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-840,-3622.5,-840,-3616.5</points>
<connection>
<GID>2282</GID>
<name>IN_1</name></connection>
<intersection>-3616.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-840,-3616.5,-829,-3616.5</points>
<intersection>-840 1</intersection>
<intersection>-829 0</intersection></hsegment></shape></wire>
<wire>
<ID>2411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-817.5,-3617.5,-817.5,-3610.5</points>
<connection>
<GID>2261</GID>
<name>OUT_0</name></connection>
<intersection>-3617.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-838,-3622.5,-838,-3617.5</points>
<connection>
<GID>2282</GID>
<name>IN_0</name></connection>
<intersection>-3617.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-838,-3617.5,-817.5,-3617.5</points>
<intersection>-838 1</intersection>
<intersection>-817.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-804.5,-3616,-804.5,-3611</points>
<connection>
<GID>2263</GID>
<name>OUT_0</name></connection>
<intersection>-3616 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-805.5,-3621.5,-805.5,-3616</points>
<connection>
<GID>2293</GID>
<name>IN_1</name></connection>
<intersection>-3616 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-805.5,-3616,-804.5,-3616</points>
<intersection>-805.5 1</intersection>
<intersection>-804.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-791.5,-3616,-791.5,-3610.5</points>
<connection>
<GID>2266</GID>
<name>OUT_0</name></connection>
<intersection>-3616 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-803.5,-3621.5,-803.5,-3616</points>
<connection>
<GID>2293</GID>
<name>IN_0</name></connection>
<intersection>-3616 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-803.5,-3616,-791.5,-3616</points>
<intersection>-803.5 1</intersection>
<intersection>-791.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-841,-3632,-841,-3628.5</points>
<connection>
<GID>2282</GID>
<name>OUT</name></connection>
<intersection>-3632 9</intersection>
<intersection>-3631.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-828,-3644.5,-828,-3631.5</points>
<connection>
<GID>2296</GID>
<name>IN_1</name></connection>
<intersection>-3639.5 7</intersection>
<intersection>-3631.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-841,-3631.5,-828,-3631.5</points>
<intersection>-841 0</intersection>
<intersection>-828 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-828,-3639.5,-816.5,-3639.5</points>
<connection>
<GID>1961</GID>
<name>IN_0</name></connection>
<intersection>-828 1</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-938,-3632,-841,-3632</points>
<connection>
<GID>2047</GID>
<name>IN_0</name></connection>
<intersection>-841 0</intersection></hsegment></shape></wire>
<wire>
<ID>2415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-804.5,-3631,-804.5,-3627.5</points>
<connection>
<GID>2293</GID>
<name>OUT</name></connection>
<intersection>-3631 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-826,-3644.5,-826,-3631</points>
<connection>
<GID>2296</GID>
<name>IN_0</name></connection>
<intersection>-3641.5 6</intersection>
<intersection>-3636 7</intersection>
<intersection>-3631 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-826,-3631,-804.5,-3631</points>
<intersection>-826 1</intersection>
<intersection>-804.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-826,-3641.5,-816.5,-3641.5</points>
<connection>
<GID>1961</GID>
<name>IN_1</name></connection>
<intersection>-826 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-949,-3636,-826,-3636</points>
<connection>
<GID>2037</GID>
<name>IN_0</name></connection>
<intersection>-826 1</intersection></hsegment></shape></wire>
<wire>
<ID>2416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-822.5,-4497,-822.5,-4489.5</points>
<connection>
<GID>2172</GID>
<name>IN_0</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-825.5,-4489.5,-822.5,-4489.5</points>
<connection>
<GID>2155</GID>
<name>OUT_0</name></connection>
<intersection>-822.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-807.5,-4497,-807.5,-4489.5</points>
<connection>
<GID>2173</GID>
<name>IN_0</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-811.5,-4489.5,-807.5,-4489.5</points>
<connection>
<GID>2156</GID>
<name>OUT_0</name></connection>
<intersection>-807.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-796,-4496.5,-796,-4489.5</points>
<connection>
<GID>2176</GID>
<name>IN_0</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-797,-4489.5,-796,-4489.5</points>
<connection>
<GID>2157</GID>
<name>OUT_0</name></connection>
<intersection>-796 0</intersection></hsegment></shape></wire>
<wire>
<ID>2419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1425,-3370.5,-1417.5,-3370.5</points>
<connection>
<GID>2330</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2329</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1375.5,-3372.5,-1367.5,-3372.5</points>
<connection>
<GID>2183</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2341</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1371.5,-3381,-1371.5,-3375.5</points>
<intersection>-3381 2</intersection>
<intersection>-3375.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1371.5,-3375.5,-1367.5,-3375.5</points>
<connection>
<GID>2341</GID>
<name>clock</name></connection>
<intersection>-1371.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1417.5,-3381,-1371.5,-3381</points>
<intersection>-1417.5 3</intersection>
<intersection>-1375.5 4</intersection>
<intersection>-1371.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1417.5,-3381,-1417.5,-3373.5</points>
<connection>
<GID>2329</GID>
<name>clock</name></connection>
<intersection>-3381 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1375.5,-3381,-1375.5,-3378</points>
<connection>
<GID>2342</GID>
<name>CLK</name></connection>
<intersection>-3381 2</intersection></vsegment></shape></wire>
<wire>
<ID>2422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1397,-3384.5,-1397,-3364.5</points>
<connection>
<GID>2333</GID>
<name>IN_1</name></connection>
<intersection>-3384.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1397,-3384.5,-1361.5,-3384.5</points>
<intersection>-1397 0</intersection>
<intersection>-1361.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-1361.5,-3384.5,-1361.5,-3375.5</points>
<connection>
<GID>2341</GID>
<name>OUTINV_0</name></connection>
<intersection>-3384.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1399,-3370.5,-1399,-3364.5</points>
<connection>
<GID>2333</GID>
<name>IN_0</name></connection>
<intersection>-3370.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1411.5,-3370.5,-1399,-3370.5</points>
<connection>
<GID>2329</GID>
<name>OUT_0</name></connection>
<intersection>-1399 0</intersection></hsegment></shape></wire>
<wire>
<ID>2424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1398,-3358.5,-1398,-3206.5</points>
<connection>
<GID>2333</GID>
<name>OUT</name></connection>
<intersection>-3206.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1398,-3206.5,-1361.5,-3206.5</points>
<connection>
<GID>2328</GID>
<name>IN_1</name></connection>
<intersection>-1398 0</intersection></hsegment></shape></wire>
<wire>
<ID>2425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1411.5,-3373.5,-1406,-3373.5</points>
<connection>
<GID>2329</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>2338</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1364.5,-3413.5,-1364.5,-3378.5</points>
<connection>
<GID>2341</GID>
<name>clear</name></connection>
<intersection>-3413.5 3</intersection>
<intersection>-3386 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1402,-3386,-1364.5,-3386</points>
<intersection>-1402 2</intersection>
<intersection>-1364.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-1402,-3386,-1402,-3373.5</points>
<connection>
<GID>2338</GID>
<name>OUT_0</name></connection>
<intersection>-3386 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-1364.5,-3413.5,-1349,-3413.5</points>
<connection>
<GID>2215</GID>
<name>clear</name></connection>
<intersection>-1364.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1060.5,-3431,-1060.5,-3375.5</points>
<intersection>-3431 2</intersection>
<intersection>-3375.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1065.5,-3375.5,-1060.5,-3375.5</points>
<connection>
<GID>2185</GID>
<name>OUT</name></connection>
<intersection>-1060.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1285.5,-3431,-1060.5,-3431</points>
<intersection>-1285.5 15</intersection>
<intersection>-1236 14</intersection>
<intersection>-1210 10</intersection>
<intersection>-1180 18</intersection>
<intersection>-1141.5 16</intersection>
<intersection>-1093 17</intersection>
<intersection>-1060.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-1210,-3431,-1210,-3405</points>
<connection>
<GID>2190</GID>
<name>clear</name></connection>
<intersection>-3431 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-1236,-3431,-1236,-3405.5</points>
<connection>
<GID>2188</GID>
<name>clear</name></connection>
<intersection>-3431 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-1285.5,-3431,-1285.5,-3405</points>
<connection>
<GID>2187</GID>
<name>clear</name></connection>
<intersection>-3431 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-1141.5,-3431,-1141.5,-3407.5</points>
<connection>
<GID>2192</GID>
<name>clear</name></connection>
<intersection>-3431 2</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-1093,-3431,-1093,-3408</points>
<connection>
<GID>2193</GID>
<name>clear</name></connection>
<intersection>-3431 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-1180,-3431,-1180,-3405.5</points>
<connection>
<GID>2191</GID>
<name>clear</name></connection>
<intersection>-3431 2</intersection></vsegment></shape></wire>
<wire>
<ID>2428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1276.5,-3443.5,-1276.5,-3393</points>
<intersection>-3443.5 8</intersection>
<intersection>-3437.5 5</intersection>
<intersection>-3428 3</intersection>
<intersection>-3399 2</intersection>
<intersection>-3393 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1276.5,-3393,-1272,-3393</points>
<connection>
<GID>2195</GID>
<name>IN_1</name></connection>
<intersection>-1276.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1282.5,-3399,-1276.5,-3399</points>
<connection>
<GID>2187</GID>
<name>Q</name></connection>
<intersection>-1276.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1276.5,-3428,-1073.5,-3428</points>
<connection>
<GID>2214</GID>
<name>IN_0</name></connection>
<intersection>-1276.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1276.5,-3437.5,-1257.5,-3437.5</points>
<intersection>-1276.5 0</intersection>
<intersection>-1257.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-1257.5,-3470,-1257.5,-3437.5</points>
<connection>
<GID>2238</GID>
<name>IN_0</name></connection>
<intersection>-3437.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1276.5,-3443.5,-1270.5,-3443.5</points>
<connection>
<GID>2186</GID>
<name>IN_0</name></connection>
<intersection>-1276.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1280.5,-3408.5,-1280.5,-3403</points>
<intersection>-3408.5 3</intersection>
<intersection>-3403 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1282.5,-3403,-1280.5,-3403</points>
<connection>
<GID>2187</GID>
<name>nQ</name></connection>
<intersection>-1280.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1280.5,-3408.5,-1273,-3408.5</points>
<connection>
<GID>2197</GID>
<name>IN_0</name></connection>
<intersection>-1280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1262,-3400.5,-1262,-3391</points>
<intersection>-3400.5 1</intersection>
<intersection>-3392 2</intersection>
<intersection>-3391 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1262,-3400.5,-1258,-3400.5</points>
<connection>
<GID>2207</GID>
<name>IN_0</name></connection>
<intersection>-1262 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1266,-3392,-1262,-3392</points>
<connection>
<GID>2195</GID>
<name>OUT</name></connection>
<intersection>-1262 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1262,-3391,-1231,-3391</points>
<connection>
<GID>2198</GID>
<name>IN_0</name></connection>
<intersection>-1262 0</intersection></hsegment></shape></wire>
<wire>
<ID>2431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1261.5,-3411.5,-1261.5,-3402.5</points>
<intersection>-3411.5 2</intersection>
<intersection>-3409.5 3</intersection>
<intersection>-3402.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1261.5,-3402.5,-1258,-3402.5</points>
<connection>
<GID>2207</GID>
<name>IN_1</name></connection>
<intersection>-1261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1261.5,-3411.5,-1228.5,-3411.5</points>
<connection>
<GID>2199</GID>
<name>IN_1</name></connection>
<intersection>-1261.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1267,-3409.5,-1261.5,-3409.5</points>
<connection>
<GID>2197</GID>
<name>OUT</name></connection>
<intersection>-1261.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1232,-3469.5,-1232,-3393</points>
<intersection>-3469.5 9</intersection>
<intersection>-3443 5</intersection>
<intersection>-3427 3</intersection>
<intersection>-3399.5 2</intersection>
<intersection>-3393 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1232,-3393,-1231,-3393</points>
<connection>
<GID>2198</GID>
<name>IN_1</name></connection>
<intersection>-1232 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1233,-3399.5,-1232,-3399.5</points>
<connection>
<GID>2188</GID>
<name>Q</name></connection>
<intersection>-1232 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1232,-3427,-1073.5,-3427</points>
<connection>
<GID>2214</GID>
<name>IN_1</name></connection>
<intersection>-1232 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1232,-3443,-1227.5,-3443</points>
<connection>
<GID>2189</GID>
<name>IN_0</name></connection>
<intersection>-1232 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1245,-3469.5,-1232,-3469.5</points>
<intersection>-1245 10</intersection>
<intersection>-1232 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-1245,-3471,-1245,-3469.5</points>
<connection>
<GID>2239</GID>
<name>IN_0</name></connection>
<intersection>-3469.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>2433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1261.5,-3711,-1261.5,-3443.5</points>
<intersection>-3711 12</intersection>
<intersection>-3555 5</intersection>
<intersection>-3458.5 10</intersection>
<intersection>-3443.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1264.5,-3443.5,-1261.5,-3443.5</points>
<connection>
<GID>2186</GID>
<name>OUT_0</name></connection>
<intersection>-1261.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1261.5,-3555,-959,-3555</points>
<intersection>-1261.5 0</intersection>
<intersection>-959 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-959,-3555,-959,-3554.5</points>
<connection>
<GID>2171</GID>
<name>IN_1</name></connection>
<intersection>-3555 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-1261.5,-3458.5,-1054,-3458.5</points>
<connection>
<GID>2217</GID>
<name>IN_0</name></connection>
<intersection>-1261.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-1261.5,-3711,-962,-3711</points>
<connection>
<GID>2346</GID>
<name>IN_1</name></connection>
<intersection>-1261.5 0</intersection>
<intersection>-1261 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-1261,-4222.5,-1261,-3711</points>
<intersection>-4222.5 19</intersection>
<intersection>-4023.5 17</intersection>
<intersection>-3841.5 15</intersection>
<intersection>-3711 12</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-1261,-3841.5,-949.5,-3841.5</points>
<connection>
<GID>1950</GID>
<name>IN_1</name></connection>
<intersection>-1261 14</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-1261,-4023.5,-941.5,-4023.5</points>
<connection>
<GID>2025</GID>
<name>IN_1</name></connection>
<intersection>-1261 14</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-1261,-4222.5,-931,-4222.5</points>
<connection>
<GID>2141</GID>
<name>IN_1</name></connection>
<intersection>-1261 14</intersection>
<intersection>-1260 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-1260,-4444.5,-1260,-4222.5</points>
<intersection>-4444.5 21</intersection>
<intersection>-4222.5 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-1260,-4444.5,-937.5,-4444.5</points>
<connection>
<GID>2394</GID>
<name>IN_1</name></connection>
<intersection>-1260 20</intersection>
<intersection>-1259 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-1259,-4678.5,-1259,-4444.5</points>
<intersection>-4678.5 23</intersection>
<intersection>-4444.5 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>-1259,-4678.5,-935.5,-4678.5</points>
<connection>
<GID>2434</GID>
<name>IN_1</name></connection>
<intersection>-1259 22</intersection>
<intersection>-1257.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-1257.5,-4905.5,-1257.5,-4678.5</points>
<intersection>-4905.5 25</intersection>
<intersection>-4678.5 23</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>-1257.5,-4905.5,-926.5,-4905.5</points>
<connection>
<GID>2472</GID>
<name>IN_1</name></connection>
<intersection>-1257.5 24</intersection></hsegment></shape></wire>
<wire>
<ID>2434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1223.5,-3392.5,-1223.5,-3392</points>
<intersection>-3392.5 2</intersection>
<intersection>-3392 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1225,-3392,-1223.5,-3392</points>
<connection>
<GID>2198</GID>
<name>OUT</name></connection>
<intersection>-1223.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1223.5,-3392.5,-1201.5,-3392.5</points>
<connection>
<GID>2200</GID>
<name>IN_0</name></connection>
<intersection>-1223.5 0</intersection>
<intersection>-1221.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-1221.5,-3399.5,-1221.5,-3392.5</points>
<connection>
<GID>2209</GID>
<name>IN_0</name></connection>
<intersection>-3392.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>2435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1230.5,-3409.5,-1230.5,-3403.5</points>
<intersection>-3409.5 2</intersection>
<intersection>-3403.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1233,-3403.5,-1230.5,-3403.5</points>
<connection>
<GID>2188</GID>
<name>nQ</name></connection>
<intersection>-1230.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1230.5,-3409.5,-1228.5,-3409.5</points>
<connection>
<GID>2199</GID>
<name>IN_0</name></connection>
<intersection>-1230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1222,-3413,-1222,-3401.5</points>
<intersection>-3413 3</intersection>
<intersection>-3410.5 1</intersection>
<intersection>-3401.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1222.5,-3410.5,-1222,-3410.5</points>
<connection>
<GID>2199</GID>
<name>OUT</name></connection>
<intersection>-1222 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1222,-3401.5,-1221.5,-3401.5</points>
<connection>
<GID>2209</GID>
<name>IN_1</name></connection>
<intersection>-1222 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1222,-3413,-1199,-3413</points>
<connection>
<GID>2201</GID>
<name>IN_1</name></connection>
<intersection>-1222 0</intersection></hsegment></shape></wire>
<wire>
<ID>2437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1205,-3470,-1205,-3372.5</points>
<intersection>-3470 13</intersection>
<intersection>-3443 9</intersection>
<intersection>-3426 2</intersection>
<intersection>-3399 1</intersection>
<intersection>-3394.5 5</intersection>
<intersection>-3372.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1207,-3399,-1205,-3399</points>
<connection>
<GID>2190</GID>
<name>Q</name></connection>
<intersection>-1205 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1205,-3426,-1073.5,-3426</points>
<connection>
<GID>2214</GID>
<name>IN_2</name></connection>
<intersection>-1205 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1205,-3394.5,-1201.5,-3394.5</points>
<connection>
<GID>2200</GID>
<name>IN_1</name></connection>
<intersection>-1205 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1205,-3372.5,-1071.5,-3372.5</points>
<connection>
<GID>2185</GID>
<name>IN_0</name></connection>
<intersection>-1205 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1205,-3443,-1198,-3443</points>
<connection>
<GID>2194</GID>
<name>IN_0</name></connection>
<intersection>-1205 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-1205,-3470,-1181,-3470</points>
<connection>
<GID>2240</GID>
<name>IN_0</name></connection>
<intersection>-1205 0</intersection></hsegment></shape></wire>
<wire>
<ID>2438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1195.5,-3393.5,-1175,-3393.5</points>
<connection>
<GID>2200</GID>
<name>OUT</name></connection>
<connection>
<GID>2202</GID>
<name>IN_0</name></connection>
<intersection>-1193 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1193,-3400,-1193,-3393.5</points>
<connection>
<GID>2210</GID>
<name>IN_0</name></connection>
<intersection>-3393.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1193,-3413,-1193,-3402</points>
<connection>
<GID>2210</GID>
<name>IN_1</name></connection>
<connection>
<GID>2201</GID>
<name>OUT</name></connection>
<intersection>-3413 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1193,-3413,-1173.5,-3413</points>
<connection>
<GID>2203</GID>
<name>IN_1</name></connection>
<intersection>-1193 0</intersection></hsegment></shape></wire>
<wire>
<ID>2440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1203.5,-3411,-1203.5,-3403</points>
<intersection>-3411 2</intersection>
<intersection>-3403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1207,-3403,-1203.5,-3403</points>
<connection>
<GID>2190</GID>
<name>nQ</name></connection>
<intersection>-1203.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1203.5,-3411,-1199,-3411</points>
<connection>
<GID>2201</GID>
<name>IN_0</name></connection>
<intersection>-1203.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1177,-3443,-1177,-3374.5</points>
<connection>
<GID>2191</GID>
<name>Q</name></connection>
<intersection>-3443 10</intersection>
<intersection>-3425 2</intersection>
<intersection>-3395.5 6</intersection>
<intersection>-3374.5 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1177,-3425,-1073.5,-3425</points>
<connection>
<GID>2214</GID>
<name>IN_3</name></connection>
<intersection>-1177 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-1177,-3395.5,-1175,-3395.5</points>
<connection>
<GID>2202</GID>
<name>IN_1</name></connection>
<intersection>-1177 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1177,-3374.5,-1071.5,-3374.5</points>
<connection>
<GID>2185</GID>
<name>IN_1</name></connection>
<intersection>-1177 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-1177,-3443,-1169.5,-3443</points>
<connection>
<GID>2206</GID>
<name>IN_0</name></connection>
<intersection>-1177 0</intersection>
<intersection>-1174 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-1174,-3470,-1174,-3443</points>
<connection>
<GID>2241</GID>
<name>IN_0</name></connection>
<intersection>-3443 10</intersection></vsegment></shape></wire>
<wire>
<ID>2442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1176,-3411,-1176,-3403.5</points>
<intersection>-3411 2</intersection>
<intersection>-3403.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1177,-3403.5,-1176,-3403.5</points>
<connection>
<GID>2191</GID>
<name>nQ</name></connection>
<intersection>-1176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1176,-3411,-1173.5,-3411</points>
<connection>
<GID>2203</GID>
<name>IN_0</name></connection>
<intersection>-1176 0</intersection></hsegment></shape></wire>
<wire>
<ID>2443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1166,-3400.5,-1166,-3392.5</points>
<intersection>-3400.5 2</intersection>
<intersection>-3394.5 1</intersection>
<intersection>-3392.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1169,-3394.5,-1166,-3394.5</points>
<connection>
<GID>2202</GID>
<name>OUT</name></connection>
<intersection>-1166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1166,-3400.5,-1164,-3400.5</points>
<connection>
<GID>2211</GID>
<name>IN_0</name></connection>
<intersection>-1166 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1166,-3392.5,-1128,-3392.5</points>
<connection>
<GID>2204</GID>
<name>IN_0</name></connection>
<intersection>-1166 0</intersection></hsegment></shape></wire>
<wire>
<ID>2444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1165.5,-3412,-1165.5,-3402.5</points>
<intersection>-3412 1</intersection>
<intersection>-3402.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1167.5,-3412,-1127.5,-3412</points>
<connection>
<GID>2203</GID>
<name>OUT</name></connection>
<connection>
<GID>2205</GID>
<name>IN_1</name></connection>
<intersection>-1165.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-1165.5,-3402.5,-1164,-3402.5</points>
<connection>
<GID>2211</GID>
<name>IN_1</name></connection>
<intersection>-1165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1133.5,-3469.5,-1133.5,-3376.5</points>
<intersection>-3469.5 14</intersection>
<intersection>-3443 9</intersection>
<intersection>-3424 3</intersection>
<intersection>-3401.5 1</intersection>
<intersection>-3394.5 10</intersection>
<intersection>-3376.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1138.5,-3401.5,-1133.5,-3401.5</points>
<connection>
<GID>2192</GID>
<name>Q</name></connection>
<intersection>-1133.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1133.5,-3424,-1073.5,-3424</points>
<connection>
<GID>2214</GID>
<name>IN_4</name></connection>
<intersection>-1133.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1133.5,-3376.5,-1071.5,-3376.5</points>
<connection>
<GID>2185</GID>
<name>IN_2</name></connection>
<intersection>-1133.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1133.5,-3443,-1123.5,-3443</points>
<connection>
<GID>2208</GID>
<name>IN_0</name></connection>
<intersection>-1133.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-1133.5,-3394.5,-1128,-3394.5</points>
<connection>
<GID>2204</GID>
<name>IN_1</name></connection>
<intersection>-1133.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-1133.5,-3469.5,-1116.5,-3469.5</points>
<connection>
<GID>2243</GID>
<name>IN_0</name></connection>
<intersection>-1133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1136,-3410,-1136,-3405.5</points>
<intersection>-3410 2</intersection>
<intersection>-3405.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1138.5,-3405.5,-1136,-3405.5</points>
<connection>
<GID>2192</GID>
<name>nQ</name></connection>
<intersection>-1136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1136,-3410,-1127.5,-3410</points>
<connection>
<GID>2205</GID>
<name>IN_0</name></connection>
<intersection>-1136 0</intersection></hsegment></shape></wire>
<wire>
<ID>2447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1121,-3401,-1121,-3393.5</points>
<intersection>-3401 2</intersection>
<intersection>-3393.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1122,-3393.5,-1121,-3393.5</points>
<connection>
<GID>2204</GID>
<name>OUT</name></connection>
<intersection>-1121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1121,-3401,-1120,-3401</points>
<connection>
<GID>2212</GID>
<name>IN_0</name></connection>
<intersection>-1121 0</intersection></hsegment></shape></wire>
<wire>
<ID>2448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1121,-3411,-1121,-3403</points>
<intersection>-3411 1</intersection>
<intersection>-3403 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1121.5,-3411,-1121,-3411</points>
<connection>
<GID>2205</GID>
<name>OUT</name></connection>
<intersection>-1121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1121,-3403,-1120,-3403</points>
<connection>
<GID>2212</GID>
<name>IN_1</name></connection>
<intersection>-1121 0</intersection></hsegment></shape></wire>
<wire>
<ID>2449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1314,-3420.5,-1096,-3420.5</points>
<intersection>-1314 16</intersection>
<intersection>-1296.5 13</intersection>
<intersection>-1239.5 12</intersection>
<intersection>-1214 6</intersection>
<intersection>-1186 7</intersection>
<intersection>-1148 11</intersection>
<intersection>-1096 28</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1214,-3420.5,-1214,-3401</points>
<intersection>-3420.5 1</intersection>
<intersection>-3401 19</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-1186,-3420.5,-1186,-3401.5</points>
<intersection>-3420.5 1</intersection>
<intersection>-3401.5 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-1148,-3420.5,-1148,-3403.5</points>
<intersection>-3420.5 1</intersection>
<intersection>-3403.5 18</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-1239.5,-3420.5,-1239.5,-3401.5</points>
<intersection>-3420.5 1</intersection>
<intersection>-3401.5 22</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-1296.5,-3420.5,-1296.5,-3401</points>
<intersection>-3420.5 1</intersection>
<intersection>-3401 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-1186,-3401.5,-1183,-3401.5</points>
<connection>
<GID>2191</GID>
<name>clock</name></connection>
<intersection>-1186 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-1296.5,-3401,-1288.5,-3401</points>
<connection>
<GID>2187</GID>
<name>clock</name></connection>
<intersection>-1296.5 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-1314,-3450,-1314,-3420.5</points>
<intersection>-3450 17</intersection>
<intersection>-3421 37</intersection>
<intersection>-3420.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-1314,-3450,-1075.5,-3450</points>
<intersection>-1314 16</intersection>
<intersection>-1270.5 34</intersection>
<intersection>-1227.5 25</intersection>
<intersection>-1198 26</intersection>
<intersection>-1169.5 24</intersection>
<intersection>-1124.5 23</intersection>
<intersection>-1075.5 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-1148,-3403.5,-1144.5,-3403.5</points>
<connection>
<GID>2192</GID>
<name>clock</name></connection>
<intersection>-1148 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-1214,-3401,-1213,-3401</points>
<connection>
<GID>2190</GID>
<name>clock</name></connection>
<intersection>-1214 6</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-1239.5,-3401.5,-1239,-3401.5</points>
<connection>
<GID>2188</GID>
<name>clock</name></connection>
<intersection>-1239.5 12</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-1124.5,-3450,-1124.5,-3446</points>
<intersection>-3450 17</intersection>
<intersection>-3446 36</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-1169.5,-3450,-1169.5,-3446</points>
<connection>
<GID>2206</GID>
<name>clock</name></connection>
<intersection>-3450 17</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>-1227.5,-3450,-1227.5,-3446</points>
<connection>
<GID>2189</GID>
<name>clock</name></connection>
<intersection>-3450 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-1198,-3450,-1198,-3446</points>
<connection>
<GID>2194</GID>
<name>clock</name></connection>
<intersection>-3450 17</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-1096,-3420.5,-1096,-3404</points>
<connection>
<GID>2193</GID>
<name>clock</name></connection>
<intersection>-3420.5 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-1270.5,-3450,-1270.5,-3446.5</points>
<connection>
<GID>2186</GID>
<name>clock</name></connection>
<intersection>-3450 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>-1075.5,-3450,-1075.5,-3446.5</points>
<connection>
<GID>2213</GID>
<name>clock</name></connection>
<intersection>-3450 17</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>-1124.5,-3446,-1123.5,-3446</points>
<connection>
<GID>2208</GID>
<name>clock</name></connection>
<intersection>-1124.5 23</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-1355,-3421,-1314,-3421</points>
<connection>
<GID>2220</GID>
<name>OUT</name></connection>
<intersection>-1352.5 38</intersection>
<intersection>-1314 16</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>-1352.5,-3421,-1352.5,-3410.5</points>
<intersection>-3421 37</intersection>
<intersection>-3410.5 39</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-1352.5,-3410.5,-1352,-3410.5</points>
<connection>
<GID>2215</GID>
<name>clock</name></connection>
<intersection>-1352.5 38</intersection></hsegment></shape></wire>
<wire>
<ID>2450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1081,-3469,-1081,-3378.5</points>
<intersection>-3469 9</intersection>
<intersection>-3443.5 13</intersection>
<intersection>-3423 2</intersection>
<intersection>-3402 11</intersection>
<intersection>-3378.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1081,-3423,-1073.5,-3423</points>
<connection>
<GID>2214</GID>
<name>IN_5</name></connection>
<intersection>-1081 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1081,-3378.5,-1071.5,-3378.5</points>
<connection>
<GID>2185</GID>
<name>IN_3</name></connection>
<intersection>-1081 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1111,-3469,-1081,-3469</points>
<connection>
<GID>2244</GID>
<name>IN_0</name></connection>
<intersection>-1081 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-1090,-3402,-1081,-3402</points>
<connection>
<GID>2193</GID>
<name>Q</name></connection>
<intersection>-1081 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-1081,-3443.5,-1075.5,-3443.5</points>
<connection>
<GID>2213</GID>
<name>IN_0</name></connection>
<intersection>-1081 0</intersection></hsegment></shape></wire>
<wire>
<ID>2451</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-1220,-4013.5,-1220,-3443</points>
<intersection>-4013.5 20</intersection>
<intersection>-3831.5 18</intersection>
<intersection>-3702.5 16</intersection>
<intersection>-3544.5 11</intersection>
<intersection>-3457.5 14</intersection>
<intersection>-3443 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1221.5,-3443,-1220,-3443</points>
<connection>
<GID>2189</GID>
<name>OUT_0</name></connection>
<intersection>-1220 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-1220,-3544.5,-959.5,-3544.5</points>
<connection>
<GID>2174</GID>
<name>IN_1</name></connection>
<intersection>-1220 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-1220,-3457.5,-1054,-3457.5</points>
<connection>
<GID>2217</GID>
<name>IN_1</name></connection>
<intersection>-1220 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-1220,-3702.5,-962.5,-3702.5</points>
<connection>
<GID>2347</GID>
<name>IN_1</name></connection>
<intersection>-1220 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-1220,-3831.5,-950,-3831.5</points>
<connection>
<GID>1951</GID>
<name>IN_1</name></connection>
<intersection>-1220 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-1220,-4013.5,-942,-4013.5</points>
<connection>
<GID>2026</GID>
<name>IN_1</name></connection>
<intersection>-1220 3</intersection>
<intersection>-1219.5 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>-1219.5,-4212.5,-1219.5,-4013.5</points>
<intersection>-4212.5 22</intersection>
<intersection>-4013.5 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>-1221.5,-4212.5,-931.5,-4212.5</points>
<connection>
<GID>2143</GID>
<name>IN_1</name></connection>
<intersection>-1221.5 23</intersection>
<intersection>-1219.5 21</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-1221.5,-4895.5,-1221.5,-4212.5</points>
<intersection>-4895.5 28</intersection>
<intersection>-4668.5 26</intersection>
<intersection>-4434.5 24</intersection>
<intersection>-4212.5 22</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-1221.5,-4434.5,-938,-4434.5</points>
<connection>
<GID>2396</GID>
<name>IN_1</name></connection>
<intersection>-1221.5 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-1221.5,-4668.5,-936,-4668.5</points>
<connection>
<GID>2435</GID>
<name>IN_1</name></connection>
<intersection>-1221.5 23</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-1221.5,-4895.5,-927,-4895.5</points>
<connection>
<GID>2473</GID>
<name>IN_1</name></connection>
<intersection>-1221.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>2452</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-1190.5,-3694,-1190.5,-3443</points>
<intersection>-3694 14</intersection>
<intersection>-3533.5 7</intersection>
<intersection>-3456.5 12</intersection>
<intersection>-3443 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1192,-3443,-1190.5,-3443</points>
<connection>
<GID>2194</GID>
<name>OUT_0</name></connection>
<intersection>-1190.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1190.5,-3533.5,-961,-3533.5</points>
<connection>
<GID>2175</GID>
<name>IN_1</name></connection>
<intersection>-1190.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-1190.5,-3456.5,-1054,-3456.5</points>
<connection>
<GID>2217</GID>
<name>IN_2</name></connection>
<intersection>-1190.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-1190.5,-3694,-963,-3694</points>
<connection>
<GID>2348</GID>
<name>IN_1</name></connection>
<intersection>-1190.5 3</intersection>
<intersection>-1190 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-1190,-4002.5,-1190,-3694</points>
<intersection>-4002.5 18</intersection>
<intersection>-3820.5 16</intersection>
<intersection>-3694 14</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-1190,-3820.5,-951.5,-3820.5</points>
<connection>
<GID>1952</GID>
<name>IN_1</name></connection>
<intersection>-1190 15</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-1190,-4002.5,-943.5,-4002.5</points>
<connection>
<GID>2027</GID>
<name>IN_1</name></connection>
<intersection>-1190 15</intersection>
<intersection>-1189.5 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-1189.5,-4201.5,-1189.5,-4002.5</points>
<intersection>-4201.5 20</intersection>
<intersection>-4002.5 18</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-1189.5,-4201.5,-933,-4201.5</points>
<connection>
<GID>2145</GID>
<name>IN_1</name></connection>
<intersection>-1189.5 19</intersection>
<intersection>-1189 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>-1189,-4423.5,-1189,-4201.5</points>
<intersection>-4423.5 22</intersection>
<intersection>-4201.5 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>-1189.5,-4423.5,-939.5,-4423.5</points>
<connection>
<GID>2397</GID>
<name>IN_1</name></connection>
<intersection>-1189.5 23</intersection>
<intersection>-1189 21</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-1189.5,-4884.5,-1189.5,-4423.5</points>
<intersection>-4884.5 26</intersection>
<intersection>-4657.5 24</intersection>
<intersection>-4423.5 22</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-1189.5,-4657.5,-937.5,-4657.5</points>
<connection>
<GID>2436</GID>
<name>IN_1</name></connection>
<intersection>-1189.5 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-1189.5,-4884.5,-928.5,-4884.5</points>
<connection>
<GID>2474</GID>
<name>IN_1</name></connection>
<intersection>-1189.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>2453</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-1163.5,-3811.5,-1163.5,-3443</points>
<connection>
<GID>2206</GID>
<name>OUT_0</name></connection>
<intersection>-3811.5 19</intersection>
<intersection>-3686 17</intersection>
<intersection>-3524.5 7</intersection>
<intersection>-3455.5 15</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1163.5,-3524.5,-961.5,-3524.5</points>
<connection>
<GID>2177</GID>
<name>IN_1</name></connection>
<intersection>-1163.5 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-1163.5,-3455.5,-1054,-3455.5</points>
<connection>
<GID>2217</GID>
<name>IN_3</name></connection>
<intersection>-1163.5 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-1163.5,-3686,-963.5,-3686</points>
<connection>
<GID>2349</GID>
<name>IN_1</name></connection>
<intersection>-1163.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-1163.5,-3811.5,-952,-3811.5</points>
<connection>
<GID>1953</GID>
<name>IN_1</name></connection>
<intersection>-1163.5 3</intersection>
<intersection>-1163 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-1163,-4414.5,-1163,-3811.5</points>
<intersection>-4414.5 25</intersection>
<intersection>-4192.5 23</intersection>
<intersection>-3993.5 21</intersection>
<intersection>-3811.5 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-1163,-3993.5,-944,-3993.5</points>
<connection>
<GID>2028</GID>
<name>IN_1</name></connection>
<intersection>-1163 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-1163,-4192.5,-933.5,-4192.5</points>
<connection>
<GID>2147</GID>
<name>IN_1</name></connection>
<intersection>-1163 20</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-1163,-4414.5,-940,-4414.5</points>
<connection>
<GID>2398</GID>
<name>IN_1</name></connection>
<intersection>-1163 20</intersection>
<intersection>-1162.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>-1162.5,-4648.5,-1162.5,-4414.5</points>
<intersection>-4648.5 27</intersection>
<intersection>-4414.5 25</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-1163,-4648.5,-938,-4648.5</points>
<connection>
<GID>2437</GID>
<name>IN_1</name></connection>
<intersection>-1163 28</intersection>
<intersection>-1162.5 26</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-1163,-4875.5,-1163,-4648.5</points>
<intersection>-4875.5 29</intersection>
<intersection>-4648.5 27</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>-1163,-4875.5,-929,-4875.5</points>
<connection>
<GID>2475</GID>
<name>IN_1</name></connection>
<intersection>-1163 28</intersection></hsegment></shape></wire>
<wire>
<ID>2454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1105.5,-3804,-1105.5,-3443</points>
<intersection>-3804 14</intersection>
<intersection>-3677.5 12</intersection>
<intersection>-3517 5</intersection>
<intersection>-3454.5 10</intersection>
<intersection>-3443 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1117.5,-3443,-1105.5,-3443</points>
<connection>
<GID>2208</GID>
<name>OUT_0</name></connection>
<intersection>-1105.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1105.5,-3517,-962.5,-3517</points>
<connection>
<GID>2180</GID>
<name>IN_1</name></connection>
<intersection>-1105.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-1105.5,-3454.5,-1054,-3454.5</points>
<connection>
<GID>2217</GID>
<name>IN_4</name></connection>
<intersection>-1105.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-1105.5,-3677.5,-964,-3677.5</points>
<connection>
<GID>2350</GID>
<name>IN_1</name></connection>
<intersection>-1105.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-1105.5,-3804,-953,-3804</points>
<connection>
<GID>1954</GID>
<name>IN_1</name></connection>
<intersection>-1105.5 0</intersection>
<intersection>-1105 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-1105,-3986,-1105,-3804</points>
<intersection>-3986 16</intersection>
<intersection>-3804 14</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-1105,-3986,-945,-3986</points>
<connection>
<GID>2039</GID>
<name>IN_1</name></connection>
<intersection>-1105 15</intersection>
<intersection>-1104.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-1104.5,-4641,-1104.5,-3986</points>
<intersection>-4641 22</intersection>
<intersection>-4407 20</intersection>
<intersection>-4185 18</intersection>
<intersection>-3986 16</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-1104.5,-4185,-934.5,-4185</points>
<connection>
<GID>2149</GID>
<name>IN_1</name></connection>
<intersection>-1104.5 17</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-1104.5,-4407,-941,-4407</points>
<connection>
<GID>2399</GID>
<name>IN_1</name></connection>
<intersection>-1104.5 17</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-1104.5,-4641,-939,-4641</points>
<connection>
<GID>2438</GID>
<name>IN_1</name></connection>
<intersection>-1104.5 17</intersection>
<intersection>-1104 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-1104,-4868,-1104,-4641</points>
<intersection>-4868 24</intersection>
<intersection>-4641 22</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-1104,-4868,-930,-4868</points>
<connection>
<GID>2476</GID>
<name>IN_1</name></connection>
<intersection>-1104 23</intersection></hsegment></shape></wire>
<wire>
<ID>2455</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-1062.5,-3669,-1062.5,-3443.5</points>
<intersection>-3669 18</intersection>
<intersection>-3509.5 10</intersection>
<intersection>-3453.5 16</intersection>
<intersection>-3443.5 13</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-1062.5,-3509.5,-963.5,-3509.5</points>
<connection>
<GID>2181</GID>
<name>IN_1</name></connection>
<intersection>-1062.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-1069.5,-3443.5,-1062.5,-3443.5</points>
<connection>
<GID>2213</GID>
<name>OUT_0</name></connection>
<intersection>-1062.5 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-1062.5,-3453.5,-1054,-3453.5</points>
<connection>
<GID>2217</GID>
<name>IN_5</name></connection>
<intersection>-1062.5 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-1062.5,-3669,-964,-3669</points>
<connection>
<GID>2351</GID>
<name>IN_1</name></connection>
<intersection>-1062.5 3</intersection>
<intersection>-1062 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-1062,-4399.5,-1062,-3669</points>
<intersection>-4399.5 26</intersection>
<intersection>-4177.5 24</intersection>
<intersection>-3978.5 22</intersection>
<intersection>-3796.5 20</intersection>
<intersection>-3669 18</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-1062,-3796.5,-954,-3796.5</points>
<connection>
<GID>1955</GID>
<name>IN_1</name></connection>
<intersection>-1062 19</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-1062,-3978.5,-946,-3978.5</points>
<connection>
<GID>2067</GID>
<name>IN_1</name></connection>
<intersection>-1062 19</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-1062,-4177.5,-935.5,-4177.5</points>
<connection>
<GID>2151</GID>
<name>IN_1</name></connection>
<intersection>-1062 19</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-1062,-4399.5,-942,-4399.5</points>
<connection>
<GID>2400</GID>
<name>IN_1</name></connection>
<intersection>-1062 19</intersection>
<intersection>-1061.5 27</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>-1061.5,-4860.5,-1061.5,-4399.5</points>
<intersection>-4860.5 30</intersection>
<intersection>-4633.5 28</intersection>
<intersection>-4399.5 26</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-1061.5,-4633.5,-940,-4633.5</points>
<connection>
<GID>2439</GID>
<name>IN_1</name></connection>
<intersection>-1061.5 27</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-1061.5,-4860.5,-931,-4860.5</points>
<connection>
<GID>2477</GID>
<name>IN_1</name></connection>
<intersection>-1061.5 27</intersection></hsegment></shape></wire>
<wire>
<ID>2456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1291.5,-3399,-1291.5,-3386.5</points>
<intersection>-3399 8</intersection>
<intersection>-3386.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-1300,-3386.5,-1291.5,-3386.5</points>
<intersection>-1300 9</intersection>
<intersection>-1291.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1291.5,-3399,-1288.5,-3399</points>
<connection>
<GID>2187</GID>
<name>J</name></connection>
<intersection>-1291.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-1300,-3387,-1300,-3375</points>
<connection>
<GID>2229</GID>
<name>IN_0</name></connection>
<intersection>-3386.5 6</intersection>
<intersection>-3375 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-1341,-3375,-1300,-3375</points>
<intersection>-1341 14</intersection>
<intersection>-1300 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-1341,-3378.5,-1341,-3375</points>
<intersection>-3378.5 15</intersection>
<intersection>-3375 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-1351.5,-3378.5,-1341,-3378.5</points>
<connection>
<GID>2247</GID>
<name>OUT</name></connection>
<intersection>-1341 14</intersection></hsegment></shape></wire>
<wire>
<ID>2457</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-1306.5,-3379.5,-1108.5,-3379.5</points>
<intersection>-1306.5 7</intersection>
<intersection>-1251 6</intersection>
<intersection>-1214.5 10</intersection>
<intersection>-1186 12</intersection>
<intersection>-1156 14</intersection>
<intersection>-1108.5 16</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1251,-3384.5,-1251,-3379.5</points>
<connection>
<GID>2231</GID>
<name>IN_1</name></connection>
<intersection>-3379.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-1306.5,-3386.5,-1306.5,-3379.5</points>
<intersection>-3386.5 20</intersection>
<intersection>-3379.5 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-1214.5,-3384,-1214.5,-3379.5</points>
<connection>
<GID>2232</GID>
<name>IN_1</name></connection>
<intersection>-3379.5 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-1186,-3384.5,-1186,-3379.5</points>
<connection>
<GID>2233</GID>
<name>IN_1</name></connection>
<intersection>-3379.5 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-1156,-3384.5,-1156,-3379.5</points>
<connection>
<GID>2234</GID>
<name>IN_1</name></connection>
<intersection>-3379.5 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-1108.5,-3382.5,-1108.5,-3379.5</points>
<connection>
<GID>2235</GID>
<name>IN_1</name></connection>
<intersection>-3379.5 4</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-1337,-3386.5,-1302,-3386.5</points>
<intersection>-1337 23</intersection>
<intersection>-1306.5 7</intersection>
<intersection>-1302 26</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-1337,-3522,-1337,-3386.5</points>
<intersection>-3522 24</intersection>
<intersection>-3386.5 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-1337,-3522,-1273,-3522</points>
<intersection>-1337 23</intersection>
<intersection>-1273 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-1273,-3522,-1273,-3521</points>
<connection>
<GID>2236</GID>
<name>OUT</name></connection>
<intersection>-3522 24</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-1302,-3387,-1302,-3386.5</points>
<connection>
<GID>2229</GID>
<name>IN_1</name></connection>
<intersection>-3386.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>2458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1301,-3403,-1301,-3393</points>
<connection>
<GID>2229</GID>
<name>OUT</name></connection>
<intersection>-3403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1301,-3403,-1288.5,-3403</points>
<connection>
<GID>2187</GID>
<name>K</name></connection>
<intersection>-1301 0</intersection></hsegment></shape></wire>
<wire>
<ID>2459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1252.5,-3493,-1252.5,-3481.5</points>
<connection>
<GID>2223</GID>
<name>IN_1</name></connection>
<intersection>-3481.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1257.5,-3481.5,-1257.5,-3476</points>
<connection>
<GID>2238</GID>
<name>OUT_0</name></connection>
<intersection>-3481.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1257.5,-3481.5,-1252.5,-3481.5</points>
<intersection>-1257.5 1</intersection>
<intersection>-1252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1250.5,-3493,-1250.5,-3481.5</points>
<connection>
<GID>2223</GID>
<name>IN_0</name></connection>
<intersection>-3481.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1245,-3481.5,-1245,-3477</points>
<connection>
<GID>2239</GID>
<name>OUT_0</name></connection>
<intersection>-3481.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1250.5,-3481.5,-1245,-3481.5</points>
<intersection>-1250.5 0</intersection>
<intersection>-1245 1</intersection></hsegment></shape></wire>
<wire>
<ID>2461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1274,-3515,-1274,-3502.5</points>
<connection>
<GID>2236</GID>
<name>IN_2</name></connection>
<intersection>-3502.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1251.5,-3502.5,-1251.5,-3499</points>
<connection>
<GID>2223</GID>
<name>OUT</name></connection>
<intersection>-3502.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1274,-3502.5,-1251.5,-3502.5</points>
<intersection>-1274 0</intersection>
<intersection>-1251.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1176.5,-3479.5,-1176.5,-3477.5</points>
<connection>
<GID>2226</GID>
<name>IN_0</name></connection>
<intersection>-3477.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1174,-3477.5,-1174,-3476</points>
<connection>
<GID>2241</GID>
<name>OUT_0</name></connection>
<intersection>-3477.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1176.5,-3477.5,-1174,-3477.5</points>
<intersection>-1176.5 0</intersection>
<intersection>-1174 1</intersection></hsegment></shape></wire>
<wire>
<ID>2463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1178.5,-3479.5,-1178.5,-3477.5</points>
<connection>
<GID>2226</GID>
<name>IN_1</name></connection>
<intersection>-3477.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1181,-3477.5,-1181,-3476</points>
<connection>
<GID>2240</GID>
<name>OUT_0</name></connection>
<intersection>-3477.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1181,-3477.5,-1178.5,-3477.5</points>
<intersection>-1181 1</intersection>
<intersection>-1178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1272,-3515,-1272,-3504.5</points>
<connection>
<GID>2236</GID>
<name>IN_1</name></connection>
<intersection>-3504.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1177.5,-3504.5,-1177.5,-3485.5</points>
<connection>
<GID>2226</GID>
<name>OUT</name></connection>
<intersection>-3504.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1272,-3504.5,-1177.5,-3504.5</points>
<intersection>-1272 0</intersection>
<intersection>-1177.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1113.5,-3478,-1113.5,-3476.5</points>
<connection>
<GID>2228</GID>
<name>IN_0</name></connection>
<intersection>-3476.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1111,-3476.5,-1111,-3475</points>
<connection>
<GID>2244</GID>
<name>OUT_0</name></connection>
<intersection>-3476.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1113.5,-3476.5,-1111,-3476.5</points>
<intersection>-1113.5 0</intersection>
<intersection>-1111 1</intersection></hsegment></shape></wire>
<wire>
<ID>2466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1115.5,-3478,-1115.5,-3476.5</points>
<connection>
<GID>2228</GID>
<name>IN_1</name></connection>
<intersection>-3476.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1116.5,-3476.5,-1116.5,-3475.5</points>
<connection>
<GID>2243</GID>
<name>OUT_0</name></connection>
<intersection>-3476.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1116.5,-3476.5,-1115.5,-3476.5</points>
<intersection>-1116.5 1</intersection>
<intersection>-1115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1270,-3515,-1270,-3507</points>
<connection>
<GID>2236</GID>
<name>IN_0</name></connection>
<intersection>-3507 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1114.5,-3507,-1114.5,-3484</points>
<connection>
<GID>2228</GID>
<name>OUT</name></connection>
<intersection>-3507 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1270,-3507,-1114.5,-3507</points>
<intersection>-1270 0</intersection>
<intersection>-1114.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1241.5,-3401.5,-1241.5,-3384</points>
<intersection>-3401.5 2</intersection>
<intersection>-3399.5 1</intersection>
<intersection>-3384 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1241.5,-3399.5,-1239,-3399.5</points>
<connection>
<GID>2188</GID>
<name>J</name></connection>
<intersection>-1241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1252,-3401.5,-1241.5,-3401.5</points>
<connection>
<GID>2207</GID>
<name>OUT</name></connection>
<intersection>-1241.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1249,-3384,-1241.5,-3384</points>
<intersection>-1249 4</intersection>
<intersection>-1241.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1249,-3384.5,-1249,-3384</points>
<connection>
<GID>2231</GID>
<name>IN_0</name></connection>
<intersection>-3384 3</intersection></vsegment></shape></wire>
<wire>
<ID>2469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1250,-3403.5,-1250,-3390.5</points>
<connection>
<GID>2231</GID>
<name>OUT</name></connection>
<intersection>-3403.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1250,-3403.5,-1239,-3403.5</points>
<connection>
<GID>2188</GID>
<name>K</name></connection>
<intersection>-1250 0</intersection></hsegment></shape></wire>
<wire>
<ID>2470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1213.5,-3399,-1213.5,-3390</points>
<connection>
<GID>2232</GID>
<name>OUT</name></connection>
<intersection>-3399 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1213.5,-3399,-1213,-3399</points>
<connection>
<GID>2190</GID>
<name>J</name></connection>
<intersection>-1213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1206,-3391.5,-1206,-3384</points>
<intersection>-3391.5 1</intersection>
<intersection>-3384 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1215.5,-3391.5,-1206,-3391.5</points>
<intersection>-1215.5 4</intersection>
<intersection>-1206 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1212.5,-3384,-1206,-3384</points>
<connection>
<GID>2232</GID>
<name>IN_0</name></connection>
<intersection>-1206 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1215.5,-3403,-1215.5,-3391.5</points>
<connection>
<GID>2209</GID>
<name>OUT</name></connection>
<intersection>-3403 6</intersection>
<intersection>-3391.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-1215.5,-3403,-1213,-3403</points>
<connection>
<GID>2190</GID>
<name>K</name></connection>
<intersection>-1215.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1187,-3392,-1180.5,-3392</points>
<intersection>-1187 3</intersection>
<intersection>-1180.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1187,-3401,-1187,-3392</points>
<connection>
<GID>2210</GID>
<name>OUT</name></connection>
<intersection>-3399.5 7</intersection>
<intersection>-3392 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1180.5,-3392,-1180.5,-3384.5</points>
<intersection>-3392 1</intersection>
<intersection>-3384.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-1184,-3384.5,-1180.5,-3384.5</points>
<connection>
<GID>2233</GID>
<name>IN_0</name></connection>
<intersection>-1180.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1187,-3399.5,-1183,-3399.5</points>
<connection>
<GID>2191</GID>
<name>J</name></connection>
<intersection>-1187 3</intersection></hsegment></shape></wire>
<wire>
<ID>2473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1185,-3403.5,-1185,-3390.5</points>
<connection>
<GID>2233</GID>
<name>OUT</name></connection>
<intersection>-3403.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1185,-3403.5,-1183,-3403.5</points>
<connection>
<GID>2191</GID>
<name>K</name></connection>
<intersection>-1185 0</intersection></hsegment></shape></wire>
<wire>
<ID>2474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1158,-3401.5,-1144.5,-3401.5</points>
<connection>
<GID>2211</GID>
<name>OUT</name></connection>
<connection>
<GID>2192</GID>
<name>J</name></connection>
<intersection>-1145.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1145.5,-3401.5,-1145.5,-3383.5</points>
<intersection>-3401.5 1</intersection>
<intersection>-3383.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-1154,-3383.5,-1145.5,-3383.5</points>
<intersection>-1154 6</intersection>
<intersection>-1145.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1154,-3384.5,-1154,-3383.5</points>
<connection>
<GID>2234</GID>
<name>IN_0</name></connection>
<intersection>-3383.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>2475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1155,-3405.5,-1155,-3390.5</points>
<connection>
<GID>2234</GID>
<name>OUT</name></connection>
<intersection>-3405.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1155,-3405.5,-1144.5,-3405.5</points>
<connection>
<GID>2192</GID>
<name>K</name></connection>
<intersection>-1155 0</intersection></hsegment></shape></wire>
<wire>
<ID>2476</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1114,-3402,-1096,-3402</points>
<connection>
<GID>2212</GID>
<name>OUT</name></connection>
<connection>
<GID>2193</GID>
<name>J</name></connection>
<intersection>-1100 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1100,-3402,-1100,-3381</points>
<intersection>-3402 1</intersection>
<intersection>-3381 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1106.5,-3381,-1100,-3381</points>
<intersection>-1106.5 15</intersection>
<intersection>-1100 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-1106.5,-3382.5,-1106.5,-3381</points>
<connection>
<GID>2235</GID>
<name>IN_0</name></connection>
<intersection>-3381 8</intersection></vsegment></shape></wire>
<wire>
<ID>2477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1107.5,-3406,-1107.5,-3388.5</points>
<connection>
<GID>2235</GID>
<name>OUT</name></connection>
<intersection>-3406 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1107.5,-3406,-1096,-3406</points>
<connection>
<GID>2193</GID>
<name>K</name></connection>
<intersection>-1107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1361.5,-3372.5,-1352.5,-3372.5</points>
<connection>
<GID>2247</GID>
<name>IN_1</name></connection>
<connection>
<GID>2341</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1350.5,-3372.5,-1350.5,-3371.5</points>
<connection>
<GID>2247</GID>
<name>IN_0</name></connection>
<intersection>-3371.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1344.5,-3371.5,-1344.5,-3370</points>
<connection>
<GID>2219</GID>
<name>OUT_0</name></connection>
<intersection>-3371.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1350.5,-3371.5,-1344.5,-3371.5</points>
<intersection>-1350.5 0</intersection>
<intersection>-1344.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1365.5,-3422,-1365.5,-3397</points>
<intersection>-3422 1</intersection>
<intersection>-3397 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1393,-3422,-1361,-3422</points>
<connection>
<GID>2218</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2220</GID>
<name>IN_1</name></connection>
<intersection>-1365.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1365.5,-3397,-1360,-3397</points>
<intersection>-1365.5 0</intersection>
<intersection>-1360 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-1360,-3405.5,-1360,-3397</points>
<connection>
<GID>2224</GID>
<name>IN_0</name></connection>
<intersection>-3397 4</intersection></vsegment></shape></wire>
<wire>
<ID>2481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1379,-3420,-1379,-3404</points>
<intersection>-3420 3</intersection>
<intersection>-3404 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1394.5,-3404,-1377.5,-3404</points>
<connection>
<GID>2216</GID>
<name>OUT_0</name></connection>
<intersection>-1379 0</intersection>
<intersection>-1377.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1379,-3420,-1361,-3420</points>
<connection>
<GID>2220</GID>
<name>IN_0</name></connection>
<intersection>-1379 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1377.5,-3404.5,-1377.5,-3404</points>
<connection>
<GID>2222</GID>
<name>IN_0</name></connection>
<intersection>-3404 1</intersection></vsegment></shape></wire>
<wire>
<ID>2482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1362,-3405.5,-1362,-3404.5</points>
<connection>
<GID>2224</GID>
<name>IN_1</name></connection>
<intersection>-3404.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1373.5,-3404.5,-1362,-3404.5</points>
<connection>
<GID>2222</GID>
<name>OUT_0</name></connection>
<intersection>-1362 0</intersection></hsegment></shape></wire>
<wire>
<ID>2483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1361,-3412,-1355.5,-3412</points>
<intersection>-1361 5</intersection>
<intersection>-1355.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-1355.5,-3412,-1355.5,-3407.5</points>
<intersection>-3412 1</intersection>
<intersection>-3407.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-1361,-3412,-1361,-3411.5</points>
<connection>
<GID>2224</GID>
<name>OUT</name></connection>
<intersection>-3412 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-1355.5,-3407.5,-1352,-3407.5</points>
<connection>
<GID>2215</GID>
<name>IN_0</name></connection>
<intersection>-1355.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1341.5,-3407.5,-1341.5,-3391</points>
<intersection>-3407.5 1</intersection>
<intersection>-3391 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1346,-3407.5,-1341.5,-3407.5</points>
<connection>
<GID>2215</GID>
<name>OUT_0</name></connection>
<intersection>-1341.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1341.5,-3391,-1272,-3391</points>
<connection>
<GID>2195</GID>
<name>IN_0</name></connection>
<intersection>-1341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1346,-3410.5,-1273,-3410.5</points>
<connection>
<GID>2215</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>2197</GID>
<name>IN_1</name></connection>
<intersection>-1315.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-1315.5,-3515,-1315.5,-3410.5</points>
<intersection>-3515 8</intersection>
<intersection>-3410.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1315.5,-3515,-1276,-3515</points>
<connection>
<GID>2236</GID>
<name>IN_3</name></connection>
<intersection>-1315.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>2486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1355,-3225.5,-712,-3225.5</points>
<intersection>-1355 15</intersection>
<intersection>-1347.5 16</intersection>
<intersection>-712 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-712,-3614,-712,-3225.5</points>
<intersection>-3614 3</intersection>
<intersection>-3225.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-869,-3614,-712,-3614</points>
<intersection>-869 14</intersection>
<intersection>-853 13</intersection>
<intersection>-839.5 12</intersection>
<intersection>-824.5 11</intersection>
<intersection>-814 10</intersection>
<intersection>-801 9</intersection>
<intersection>-712 2</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-801,-3614,-801,-3602.5</points>
<connection>
<GID>2249</GID>
<name>clock</name></connection>
<intersection>-3614 3</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-814,-3614,-814,-3602.5</points>
<connection>
<GID>2242</GID>
<name>clock</name></connection>
<intersection>-3614 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-824.5,-3614,-824.5,-3602.5</points>
<connection>
<GID>2237</GID>
<name>clock</name></connection>
<intersection>-3614 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-839.5,-3614,-839.5,-3602.5</points>
<connection>
<GID>2230</GID>
<name>clock</name></connection>
<intersection>-3614 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-853,-3614,-853,-3602.5</points>
<connection>
<GID>2221</GID>
<name>clock</name></connection>
<intersection>-3614 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-869,-3657,-869,-3602</points>
<connection>
<GID>2196</GID>
<name>clock</name></connection>
<intersection>-3657 196</intersection>
<intersection>-3614 3</intersection>
<intersection>-3602 17</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-1355,-3225.5,-1355,-3215</points>
<connection>
<GID>2299</GID>
<name>CLK</name></connection>
<intersection>-3225.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-1347.5,-3225.5,-1347.5,-3215</points>
<connection>
<GID>2270</GID>
<name>IN_1</name></connection>
<intersection>-3225.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-1004.5,-3602,-869,-3602</points>
<intersection>-1004.5 18</intersection>
<intersection>-898.5 210</intersection>
<intersection>-869 14</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-1004.5,-3727,-1004.5,-3602</points>
<intersection>-3727 41</intersection>
<intersection>-3602 17</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>-1005,-3727,-802.5,-3727</points>
<connection>
<GID>2168</GID>
<name>clock</name></connection>
<intersection>-1005 89</intersection>
<intersection>-1004.5 18</intersection>
<intersection>-900 215</intersection>
<intersection>-869.5 52</intersection>
<intersection>-854 51</intersection>
<intersection>-840.5 50</intersection>
<intersection>-826.5 49</intersection>
<intersection>-815.5 48</intersection>
<intersection>-802.5 47</intersection></hsegment>
<vsegment>
<ID>47</ID>
<points>-802.5,-3727.5,-802.5,-3727</points>
<intersection>-3727.5 88</intersection>
<intersection>-3727 41</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>-815.5,-3727.5,-815.5,-3727</points>
<intersection>-3727.5 87</intersection>
<intersection>-3727 41</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>-826.5,-3727.5,-826.5,-3727</points>
<intersection>-3727.5 86</intersection>
<intersection>-3727 41</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>-840.5,-3727.5,-840.5,-3727</points>
<intersection>-3727.5 85</intersection>
<intersection>-3727 41</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>-854,-3727.5,-854,-3727</points>
<intersection>-3727.5 84</intersection>
<intersection>-3727 41</intersection></vsegment>
<vsegment>
<ID>52</ID>
<points>-869.5,-3774,-869.5,-3727</points>
<intersection>-3774 198</intersection>
<intersection>-3727 41</intersection></vsegment>
<hsegment>
<ID>84</ID>
<points>-854,-3727.5,-853.5,-3727.5</points>
<connection>
<GID>1915</GID>
<name>clock</name></connection>
<intersection>-854 51</intersection></hsegment>
<hsegment>
<ID>85</ID>
<points>-840.5,-3727.5,-840,-3727.5</points>
<connection>
<GID>1917</GID>
<name>clock</name></connection>
<intersection>-840.5 50</intersection></hsegment>
<hsegment>
<ID>86</ID>
<points>-826.5,-3727.5,-825,-3727.5</points>
<connection>
<GID>1919</GID>
<name>clock</name></connection>
<intersection>-826.5 49</intersection></hsegment>
<hsegment>
<ID>87</ID>
<points>-815.5,-3727.5,-814.5,-3727.5</points>
<connection>
<GID>1920</GID>
<name>clock</name></connection>
<intersection>-815.5 48</intersection></hsegment>
<hsegment>
<ID>88</ID>
<points>-802.5,-3727.5,-801.5,-3727.5</points>
<connection>
<GID>1921</GID>
<name>clock</name></connection>
<intersection>-802.5 47</intersection></hsegment>
<vsegment>
<ID>89</ID>
<points>-1005,-4282,-1005,-3727</points>
<intersection>-4282 109</intersection>
<intersection>-4280.5 138</intersection>
<intersection>-4070.5 122</intersection>
<intersection>-3901 93</intersection>
<intersection>-3727 41</intersection></vsegment>
<hsegment>
<ID>93</ID>
<points>-1005,-3901,-791.5,-3901</points>
<intersection>-1005 89</intersection>
<intersection>-924 213</intersection>
<intersection>-859.5 104</intersection>
<intersection>-843.5 103</intersection>
<intersection>-830 102</intersection>
<intersection>-815 101</intersection>
<intersection>-804.5 100</intersection>
<intersection>-791.5 99</intersection></hsegment>
<vsegment>
<ID>99</ID>
<points>-791.5,-3901,-791.5,-3889.5</points>
<connection>
<GID>1885</GID>
<name>clock</name></connection>
<intersection>-3901 93</intersection></vsegment>
<vsegment>
<ID>100</ID>
<points>-804.5,-3901,-804.5,-3889.5</points>
<connection>
<GID>1884</GID>
<name>clock</name></connection>
<intersection>-3901 93</intersection></vsegment>
<vsegment>
<ID>101</ID>
<points>-815,-3901,-815,-3889.5</points>
<connection>
<GID>1881</GID>
<name>clock</name></connection>
<intersection>-3901 93</intersection></vsegment>
<vsegment>
<ID>102</ID>
<points>-830,-3901,-830,-3889.5</points>
<connection>
<GID>1870</GID>
<name>clock</name></connection>
<intersection>-3901 93</intersection></vsegment>
<vsegment>
<ID>103</ID>
<points>-843.5,-3901,-843.5,-3889.5</points>
<connection>
<GID>1860</GID>
<name>clock</name></connection>
<intersection>-3901 93</intersection></vsegment>
<vsegment>
<ID>104</ID>
<points>-859.5,-3943,-859.5,-3889</points>
<connection>
<GID>1956</GID>
<name>clock</name></connection>
<intersection>-3943 200</intersection>
<intersection>-3901 93</intersection></vsegment>
<hsegment>
<ID>109</ID>
<points>-1005.5,-4282,-773,-4282</points>
<intersection>-1005.5 153</intersection>
<intersection>-1005 89</intersection>
<intersection>-909 219</intersection>
<intersection>-841 205</intersection>
<intersection>-825 119</intersection>
<intersection>-811.5 118</intersection>
<intersection>-796.5 117</intersection>
<intersection>-786 116</intersection>
<intersection>-773 115</intersection></hsegment>
<vsegment>
<ID>115</ID>
<points>-773,-4282,-773,-4270.5</points>
<connection>
<GID>2076</GID>
<name>clock</name></connection>
<intersection>-4282 109</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>-786,-4282,-786,-4270.5</points>
<connection>
<GID>2075</GID>
<name>clock</name></connection>
<intersection>-4282 109</intersection></vsegment>
<vsegment>
<ID>117</ID>
<points>-796.5,-4282,-796.5,-4270.5</points>
<connection>
<GID>2073</GID>
<name>clock</name></connection>
<intersection>-4282 109</intersection></vsegment>
<vsegment>
<ID>118</ID>
<points>-811.5,-4282,-811.5,-4270.5</points>
<connection>
<GID>2072</GID>
<name>clock</name></connection>
<intersection>-4282 109</intersection></vsegment>
<vsegment>
<ID>119</ID>
<points>-825,-4282,-825,-4270.5</points>
<connection>
<GID>2070</GID>
<name>clock</name></connection>
<intersection>-4282 109</intersection></vsegment>
<hsegment>
<ID>122</ID>
<points>-1005,-4070.5,-851.5,-4070.5</points>
<intersection>-1005 89</intersection>
<intersection>-922.5 221</intersection>
<intersection>-851.5 137</intersection></hsegment>
<hsegment>
<ID>126</ID>
<points>-851.5,-4083,-783.5,-4083</points>
<intersection>-851.5 137</intersection>
<intersection>-835.5 136</intersection>
<intersection>-822 135</intersection>
<intersection>-807 134</intersection>
<intersection>-796.5 133</intersection>
<intersection>-783.5 132</intersection></hsegment>
<vsegment>
<ID>132</ID>
<points>-783.5,-4083,-783.5,-4071.5</points>
<connection>
<GID>1997</GID>
<name>clock</name></connection>
<intersection>-4083 126</intersection></vsegment>
<vsegment>
<ID>133</ID>
<points>-796.5,-4083,-796.5,-4071.5</points>
<connection>
<GID>1996</GID>
<name>clock</name></connection>
<intersection>-4083 126</intersection></vsegment>
<vsegment>
<ID>134</ID>
<points>-807,-4083,-807,-4071.5</points>
<connection>
<GID>1995</GID>
<name>clock</name></connection>
<intersection>-4083 126</intersection></vsegment>
<vsegment>
<ID>135</ID>
<points>-822,-4083,-822,-4071.5</points>
<connection>
<GID>1994</GID>
<name>clock</name></connection>
<intersection>-4083 126</intersection></vsegment>
<vsegment>
<ID>136</ID>
<points>-835.5,-4083,-835.5,-4071.5</points>
<connection>
<GID>1993</GID>
<name>clock</name></connection>
<intersection>-4083 126</intersection></vsegment>
<vsegment>
<ID>137</ID>
<points>-851.5,-4128.5,-851.5,-4070.5</points>
<connection>
<GID>2069</GID>
<name>clock</name></connection>
<intersection>-4128.5 227</intersection>
<intersection>-4083 126</intersection>
<intersection>-4070.5 122</intersection></vsegment>
<hsegment>
<ID>138</ID>
<points>-1005.5,-4280.5,-1005,-4280.5</points>
<intersection>-1005.5 153</intersection>
<intersection>-1005 89</intersection></hsegment>
<hsegment>
<ID>142</ID>
<points>-1005.5,-4504,-779.5,-4504</points>
<intersection>-1005.5 153</intersection>
<intersection>-906 218</intersection>
<intersection>-847.5 194</intersection>
<intersection>-831.5 152</intersection>
<intersection>-818 151</intersection>
<intersection>-803 150</intersection>
<intersection>-792.5 149</intersection>
<intersection>-779.5 148</intersection></hsegment>
<vsegment>
<ID>148</ID>
<points>-779.5,-4504,-779.5,-4492.5</points>
<connection>
<GID>2169</GID>
<name>clock</name></connection>
<intersection>-4504 142</intersection></vsegment>
<vsegment>
<ID>149</ID>
<points>-792.5,-4504,-792.5,-4492.5</points>
<connection>
<GID>2158</GID>
<name>clock</name></connection>
<intersection>-4504 142</intersection></vsegment>
<vsegment>
<ID>150</ID>
<points>-803,-4504,-803,-4492.5</points>
<connection>
<GID>2157</GID>
<name>clock</name></connection>
<intersection>-4504 142</intersection></vsegment>
<vsegment>
<ID>151</ID>
<points>-818,-4504,-818,-4492.5</points>
<intersection>-4504 142</intersection>
<intersection>-4492.5 217</intersection></vsegment>
<vsegment>
<ID>152</ID>
<points>-831.5,-4504,-831.5,-4492.5</points>
<connection>
<GID>2155</GID>
<name>clock</name></connection>
<intersection>-4504 142</intersection></vsegment>
<vsegment>
<ID>153</ID>
<points>-1005.5,-4965,-1005.5,-4280.5</points>
<intersection>-4965 174</intersection>
<intersection>-4953 192</intersection>
<intersection>-4784.5 208</intersection>
<intersection>-4738 158</intersection>
<intersection>-4504 142</intersection>
<intersection>-4325 204</intersection>
<intersection>-4282 109</intersection>
<intersection>-4280.5 138</intersection></vsegment>
<hsegment>
<ID>158</ID>
<points>-1005.5,-4738,-777.5,-4738</points>
<intersection>-1005.5 153</intersection>
<intersection>-906 222</intersection>
<intersection>-845.5 169</intersection>
<intersection>-829.5 168</intersection>
<intersection>-816 167</intersection>
<intersection>-801 166</intersection>
<intersection>-790.5 209</intersection>
<intersection>-777.5 164</intersection></hsegment>
<vsegment>
<ID>164</ID>
<points>-777.5,-4738,-777.5,-4726.5</points>
<connection>
<GID>2406</GID>
<name>clock</name></connection>
<intersection>-4738 158</intersection></vsegment>
<vsegment>
<ID>166</ID>
<points>-801,-4738,-801,-4726.5</points>
<connection>
<GID>2404</GID>
<name>clock</name></connection>
<intersection>-4738 158</intersection></vsegment>
<vsegment>
<ID>167</ID>
<points>-816,-4738,-816,-4726.5</points>
<connection>
<GID>2403</GID>
<name>clock</name></connection>
<intersection>-4738 158</intersection></vsegment>
<vsegment>
<ID>168</ID>
<points>-829.5,-4738,-829.5,-4726.5</points>
<connection>
<GID>2402</GID>
<name>clock</name></connection>
<intersection>-4738 158</intersection></vsegment>
<vsegment>
<ID>169</ID>
<points>-845.5,-4738,-845.5,-4726</points>
<connection>
<GID>2440</GID>
<name>clock</name></connection>
<intersection>-4738 158</intersection></vsegment>
<hsegment>
<ID>174</ID>
<points>-1005.5,-4965,-768.5,-4965</points>
<intersection>-1005.5 153</intersection>
<intersection>-885 224</intersection>
<intersection>-820.5 184</intersection>
<intersection>-807 183</intersection>
<intersection>-792 182</intersection>
<intersection>-781.5 181</intersection>
<intersection>-768.5 180</intersection></hsegment>
<vsegment>
<ID>180</ID>
<points>-768.5,-4965,-768.5,-4953.5</points>
<connection>
<GID>2445</GID>
<name>clock</name></connection>
<intersection>-4965 174</intersection></vsegment>
<vsegment>
<ID>181</ID>
<points>-781.5,-4965,-781.5,-4953.5</points>
<connection>
<GID>2444</GID>
<name>clock</name></connection>
<intersection>-4965 174</intersection></vsegment>
<vsegment>
<ID>182</ID>
<points>-792,-4965,-792,-4953.5</points>
<connection>
<GID>2443</GID>
<name>clock</name></connection>
<intersection>-4965 174</intersection></vsegment>
<vsegment>
<ID>183</ID>
<points>-807,-4965,-807,-4953.5</points>
<connection>
<GID>2442</GID>
<name>clock</name></connection>
<intersection>-4965 174</intersection></vsegment>
<vsegment>
<ID>184</ID>
<points>-820.5,-4965,-820.5,-4953.5</points>
<connection>
<GID>2441</GID>
<name>clock</name></connection>
<intersection>-4965 174</intersection></vsegment>
<hsegment>
<ID>192</ID>
<points>-1005.5,-4953,-836.5,-4953</points>
<connection>
<GID>2478</GID>
<name>clock</name></connection>
<intersection>-1005.5 153</intersection></hsegment>
<vsegment>
<ID>194</ID>
<points>-847.5,-4550,-847.5,-4492</points>
<connection>
<GID>2401</GID>
<name>clock</name></connection>
<intersection>-4550 229</intersection>
<intersection>-4504 142</intersection></vsegment>
<hsegment>
<ID>196</ID>
<points>-869,-3657,-802,-3657</points>
<connection>
<GID>2369</GID>
<name>clock</name></connection>
<intersection>-869 14</intersection></hsegment>
<hsegment>
<ID>198</ID>
<points>-869.5,-3774,-811.5,-3774</points>
<connection>
<GID>1864</GID>
<name>clock</name></connection>
<intersection>-869.5 52</intersection></hsegment>
<hsegment>
<ID>200</ID>
<points>-859.5,-3943,-805.5,-3943</points>
<connection>
<GID>1904</GID>
<name>clock</name></connection>
<intersection>-859.5 104</intersection></hsegment>
<hsegment>
<ID>204</ID>
<points>-1005.5,-4325,-789.5,-4325</points>
<connection>
<GID>1989</GID>
<name>clock</name></connection>
<intersection>-1005.5 153</intersection></hsegment>
<vsegment>
<ID>205</ID>
<points>-841,-4282,-841,-4270</points>
<connection>
<GID>2153</GID>
<name>clock</name></connection>
<intersection>-4282 109</intersection></vsegment>
<hsegment>
<ID>208</ID>
<points>-1005.5,-4784.5,-790.5,-4784.5</points>
<connection>
<GID>2056</GID>
<name>clock</name></connection>
<intersection>-1005.5 153</intersection></hsegment>
<vsegment>
<ID>209</ID>
<points>-790.5,-4738,-790.5,-4726.5</points>
<connection>
<GID>2405</GID>
<name>clock</name></connection>
<intersection>-4738 158</intersection></vsegment>
<vsegment>
<ID>210</ID>
<points>-898.5,-3618.5,-898.5,-3602</points>
<intersection>-3618.5 211</intersection>
<intersection>-3602 17</intersection></vsegment>
<hsegment>
<ID>211</ID>
<points>-898.5,-3618.5,-894.5,-3618.5</points>
<connection>
<GID>2035</GID>
<name>clock</name></connection>
<intersection>-898.5 210</intersection></hsegment>
<vsegment>
<ID>213</ID>
<points>-924,-3914,-924,-3901</points>
<intersection>-3914 214</intersection>
<intersection>-3901 93</intersection></vsegment>
<hsegment>
<ID>214</ID>
<points>-924,-3914,-921.5,-3914</points>
<connection>
<GID>2058</GID>
<name>clock</name></connection>
<intersection>-924 213</intersection></hsegment>
<vsegment>
<ID>215</ID>
<points>-900,-3743,-900,-3727</points>
<intersection>-3743 216</intersection>
<intersection>-3727 41</intersection></vsegment>
<hsegment>
<ID>216</ID>
<points>-900,-3743,-897.5,-3743</points>
<connection>
<GID>2048</GID>
<name>clock</name></connection>
<intersection>-900 215</intersection></hsegment>
<hsegment>
<ID>217</ID>
<points>-818,-4492.5,-817.5,-4492.5</points>
<connection>
<GID>2156</GID>
<name>clock</name></connection>
<intersection>-818 151</intersection></hsegment>
<vsegment>
<ID>218</ID>
<points>-906,-4513,-906,-4504</points>
<connection>
<GID>1903</GID>
<name>clock</name></connection>
<intersection>-4504 142</intersection></vsegment>
<vsegment>
<ID>219</ID>
<points>-909,-4290,-909,-4282</points>
<intersection>-4290 220</intersection>
<intersection>-4282 109</intersection></vsegment>
<hsegment>
<ID>220</ID>
<points>-909,-4290,-904.5,-4290</points>
<connection>
<GID>1892</GID>
<name>clock</name></connection>
<intersection>-909 219</intersection></hsegment>
<vsegment>
<ID>221</ID>
<points>-922.5,-4081.5,-922.5,-4070.5</points>
<connection>
<GID>1871</GID>
<name>clock</name></connection>
<intersection>-4070.5 122</intersection></vsegment>
<vsegment>
<ID>222</ID>
<points>-906,-4746.5,-906,-4738</points>
<intersection>-4746.5 223</intersection>
<intersection>-4738 158</intersection></vsegment>
<hsegment>
<ID>223</ID>
<points>-906,-4746.5,-904,-4746.5</points>
<connection>
<GID>1963</GID>
<name>clock</name></connection>
<intersection>-906 222</intersection></hsegment>
<vsegment>
<ID>224</ID>
<points>-885,-4975,-885,-4965</points>
<intersection>-4975 225</intersection>
<intersection>-4965 174</intersection></vsegment>
<hsegment>
<ID>225</ID>
<points>-885,-4975,-881.5,-4975</points>
<connection>
<GID>1979</GID>
<name>clock</name></connection>
<intersection>-885 224</intersection></hsegment>
<hsegment>
<ID>227</ID>
<points>-851.5,-4128.5,-797.5,-4128.5</points>
<connection>
<GID>1965</GID>
<name>clock</name></connection>
<intersection>-851.5 137</intersection></hsegment>
<hsegment>
<ID>229</ID>
<points>-847.5,-4550,-795,-4550</points>
<connection>
<GID>2033</GID>
<name>clock</name></connection>
<intersection>-847.5 194</intersection></hsegment></shape></wire>
<wire>
<ID>2487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1099.5,-3278.5,-1099.5,-3277.5</points>
<intersection>-3278.5 2</intersection>
<intersection>-3277.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1104,-3277.5,-1099.5,-3277.5</points>
<connection>
<GID>2268</GID>
<name>IN_1</name></connection>
<intersection>-1099.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1099.5,-3278.5,-1094.5,-3278.5</points>
<connection>
<GID>2257</GID>
<name>Q</name></connection>
<intersection>-1099.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1330.5,-3266,-1330.5,-3261.5</points>
<intersection>-3266 1</intersection>
<intersection>-3261.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1334,-3266,-1330.5,-3266</points>
<connection>
<GID>2275</GID>
<name>IN_1</name></connection>
<intersection>-1330.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1330.5,-3261.5,-1327,-3261.5</points>
<connection>
<GID>2274</GID>
<name>OUT</name></connection>
<intersection>-1330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-783,-4497,-783,-4489.5</points>
<connection>
<GID>2178</GID>
<name>IN_0</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-786.5,-4489.5,-783,-4489.5</points>
<connection>
<GID>2158</GID>
<name>OUT_0</name></connection>
<intersection>-783 0</intersection></hsegment></shape></wire>
<wire>
<ID>2490</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1340,-3278.5,-1110,-3278.5</points>
<connection>
<GID>2300</GID>
<name>clear</name></connection>
<connection>
<GID>2288</GID>
<name>clear</name></connection>
<connection>
<GID>2290</GID>
<name>clear</name></connection>
<connection>
<GID>2292</GID>
<name>clear</name></connection>
<connection>
<GID>2298</GID>
<name>clear</name></connection>
<connection>
<GID>2268</GID>
<name>OUT</name></connection>
<intersection>-1340 6</intersection>
<intersection>-1203.5 4</intersection>
<intersection>-1158 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1158,-3279,-1158,-3278.5</points>
<connection>
<GID>2295</GID>
<name>clear</name></connection>
<intersection>-3278.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1203.5,-3314.5,-1203.5,-3278.5</points>
<intersection>-3314.5 5</intersection>
<intersection>-3278.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-1203.5,-3314.5,-1112.5,-3314.5</points>
<intersection>-1203.5 4</intersection>
<intersection>-1194.5 13</intersection>
<intersection>-1178 12</intersection>
<intersection>-1163.5 11</intersection>
<intersection>-1146.5 10</intersection>
<intersection>-1130.5 9</intersection>
<intersection>-1112.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1340,-3278.5,-1340,-3258.5</points>
<intersection>-3278.5 1</intersection>
<intersection>-3258.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1340.5,-3258.5,-1340,-3258.5</points>
<connection>
<GID>2278</GID>
<name>IN_0</name></connection>
<intersection>-1340 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-1112.5,-3314.5,-1112.5,-3313.5</points>
<connection>
<GID>2318</GID>
<name>clear</name></connection>
<intersection>-3314.5 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-1130.5,-3314.5,-1130.5,-3313.5</points>
<connection>
<GID>2317</GID>
<name>clear</name></connection>
<intersection>-3314.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-1146.5,-3314.5,-1146.5,-3313.5</points>
<connection>
<GID>2316</GID>
<name>clear</name></connection>
<intersection>-3314.5 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-1163.5,-3314.5,-1163.5,-3313.5</points>
<connection>
<GID>2314</GID>
<name>clear</name></connection>
<intersection>-3314.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-1178,-3314.5,-1178,-3313.5</points>
<connection>
<GID>2313</GID>
<name>clear</name></connection>
<intersection>-3314.5 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-1194.5,-3314.5,-1194.5,-3313.5</points>
<connection>
<GID>2311</GID>
<name>clear</name></connection>
<intersection>-3314.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>2491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1334,-3268,-1294,-3268</points>
<connection>
<GID>2275</GID>
<name>IN_0</name></connection>
<intersection>-1294 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1294,-3270,-1294,-3268</points>
<connection>
<GID>2272</GID>
<name>OUT</name></connection>
<intersection>-3268 1</intersection></vsegment></shape></wire>
<wire>
<ID>2492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1352.5,-3257.5,-1352.5,-3253.5</points>
<intersection>-3257.5 2</intersection>
<intersection>-3253.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1359,-3253.5,-1352.5,-3253.5</points>
<connection>
<GID>2280</GID>
<name>IN_1</name></connection>
<intersection>-1352.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1352.5,-3257.5,-1346.5,-3257.5</points>
<connection>
<GID>2278</GID>
<name>OUT</name></connection>
<intersection>-1352.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1106.5,-3274.5,-1106.5,-3191.5</points>
<intersection>-3274.5 2</intersection>
<intersection>-3191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1203,-3191.5,-1106.5,-3191.5</points>
<connection>
<GID>2264</GID>
<name>IN_0</name></connection>
<intersection>-1106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1106.5,-3274.5,-1094.5,-3274.5</points>
<connection>
<GID>2257</GID>
<name>nQ</name></connection>
<intersection>-1106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1332,-3205.5,-1286.5,-3205.5</points>
<connection>
<GID>2279</GID>
<name>clear</name></connection>
<connection>
<GID>2277</GID>
<name>clear</name></connection>
<connection>
<GID>2276</GID>
<name>clear</name></connection>
<intersection>-1332 13</intersection>
<intersection>-1286.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1286.5,-3206.5,-1286.5,-3205.5</points>
<connection>
<GID>2281</GID>
<name>clear</name></connection>
<intersection>-3206.5 5</intersection>
<intersection>-3205.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-1286.5,-3206.5,-1205,-3206.5</points>
<connection>
<GID>2284</GID>
<name>clear</name></connection>
<connection>
<GID>2283</GID>
<name>clear</name></connection>
<intersection>-1286.5 4</intersection>
<intersection>-1224 12</intersection>
<intersection>-1205 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-1205,-3213.5,-1205,-3206.5</points>
<connection>
<GID>2320</GID>
<name>IN_0</name></connection>
<intersection>-3206.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-1224,-3206.5,-1224,-3199.5</points>
<connection>
<GID>2285</GID>
<name>OUT</name></connection>
<intersection>-3206.5 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-1332,-3240.5,-1332,-3205.5</points>
<intersection>-3240.5 14</intersection>
<intersection>-3205.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-1332,-3240.5,-1241,-3240.5</points>
<connection>
<GID>2326</GID>
<name>clear</name></connection>
<connection>
<GID>2325</GID>
<name>clear</name></connection>
<connection>
<GID>2324</GID>
<name>clear</name></connection>
<connection>
<GID>2323</GID>
<name>clear</name></connection>
<connection>
<GID>2322</GID>
<name>clear</name></connection>
<connection>
<GID>2321</GID>
<name>clear</name></connection>
<intersection>-1332 13</intersection></hsegment></shape></wire>
<wire>
<ID>2495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1236,-3187,-1203,-3187</points>
<intersection>-1236 3</intersection>
<intersection>-1203 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1236,-3191,-1236,-3187</points>
<intersection>-3191 5</intersection>
<intersection>-3187 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1203,-3189.5,-1203,-3187</points>
<connection>
<GID>2264</GID>
<name>IN_1</name></connection>
<intersection>-3187 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-1237,-3191,-1236,-3191</points>
<connection>
<GID>2315</GID>
<name>OUT</name></connection>
<intersection>-1236 3</intersection></hsegment></shape></wire>
<wire>
<ID>2496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-770,-4496.5,-770,-4489.5</points>
<connection>
<GID>2179</GID>
<name>IN_0</name></connection>
<intersection>-4489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-773.5,-4489.5,-770,-4489.5</points>
<connection>
<GID>2169</GID>
<name>OUT_0</name></connection>
<intersection>-770 0</intersection></hsegment></shape></wire>
<wire>
<ID>2497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-837.5,-4506.5,-837.5,-4501</points>
<connection>
<GID>2170</GID>
<name>OUT_0</name></connection>
<intersection>-4506.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-822.5,-4512.5,-822.5,-4506.5</points>
<connection>
<GID>2246</GID>
<name>IN_3</name></connection>
<intersection>-4506.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-837.5,-4506.5,-822.5,-4506.5</points>
<intersection>-837.5 0</intersection>
<intersection>-822.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1351.5,-3267,-1340,-3267</points>
<connection>
<GID>2289</GID>
<name>IN_0</name></connection>
<connection>
<GID>2275</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1357.5,-3266,-1357.5,-3255.5</points>
<connection>
<GID>2289</GID>
<name>OUT</name></connection>
<intersection>-3255.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1359,-3255.5,-1357.5,-3255.5</points>
<connection>
<GID>2280</GID>
<name>IN_0</name></connection>
<intersection>-1357.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1373,-3254.5,-1365,-3254.5</points>
<connection>
<GID>2294</GID>
<name>N_in1</name></connection>
<connection>
<GID>2280</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1213.5,-3198.5,-1213.5,-3190.5</points>
<intersection>-3198.5 1</intersection>
<intersection>-3190.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1218,-3198.5,-1213.5,-3198.5</points>
<connection>
<GID>2285</GID>
<name>IN_1</name></connection>
<intersection>-1213.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1213.5,-3190.5,-1209,-3190.5</points>
<connection>
<GID>2264</GID>
<name>OUT</name></connection>
<intersection>-1213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1213.5,-3284.5,-1213.5,-3200.5</points>
<intersection>-3284.5 3</intersection>
<intersection>-3200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1218,-3200.5,-1213.5,-3200.5</points>
<connection>
<GID>2285</GID>
<name>IN_0</name></connection>
<intersection>-1213.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1355.5,-3284.5,-1104,-3284.5</points>
<connection>
<GID>2273</GID>
<name>OUT_0</name></connection>
<intersection>-1213.5 0</intersection>
<intersection>-1104 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-1104,-3284.5,-1104,-3279.5</points>
<connection>
<GID>2268</GID>
<name>IN_0</name></connection>
<intersection>-3284.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>2503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1307,-3203.5,-1307,-3191</points>
<intersection>-3203.5 4</intersection>
<intersection>-3199.5 2</intersection>
<intersection>-3191 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1308.5,-3191,-1297.5,-3191</points>
<connection>
<GID>2302</GID>
<name>OUT</name></connection>
<connection>
<GID>2306</GID>
<name>IN_0</name></connection>
<intersection>-1307 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1307,-3199.5,-1305.5,-3199.5</points>
<connection>
<GID>2279</GID>
<name>J</name></connection>
<intersection>-1307 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1307,-3203.5,-1305.5,-3203.5</points>
<connection>
<GID>2279</GID>
<name>K</name></connection>
<intersection>-1307 0</intersection></hsegment></shape></wire>
<wire>
<ID>2504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1290.5,-3204,-1290.5,-3192</points>
<intersection>-3204 4</intersection>
<intersection>-3200 2</intersection>
<intersection>-3192 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1291.5,-3192,-1282.5,-3192</points>
<connection>
<GID>2309</GID>
<name>IN_0</name></connection>
<connection>
<GID>2306</GID>
<name>OUT</name></connection>
<intersection>-1290.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1290.5,-3200,-1289.5,-3200</points>
<connection>
<GID>2281</GID>
<name>J</name></connection>
<intersection>-1290.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1290.5,-3204,-1289.5,-3204</points>
<connection>
<GID>2281</GID>
<name>K</name></connection>
<intersection>-1290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1275,-3204.5,-1275,-3193</points>
<intersection>-3204.5 4</intersection>
<intersection>-3200.5 2</intersection>
<intersection>-3193 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1276.5,-3193,-1265,-3193</points>
<connection>
<GID>2309</GID>
<name>OUT</name></connection>
<connection>
<GID>2312</GID>
<name>IN_0</name></connection>
<intersection>-1275 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1275,-3200.5,-1273.5,-3200.5</points>
<connection>
<GID>2283</GID>
<name>J</name></connection>
<intersection>-1275 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1275,-3204.5,-1273.5,-3204.5</points>
<connection>
<GID>2283</GID>
<name>K</name></connection>
<intersection>-1275 0</intersection></hsegment></shape></wire>
<wire>
<ID>2506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1258,-3204.5,-1258,-3194</points>
<intersection>-3204.5 4</intersection>
<intersection>-3200.5 2</intersection>
<intersection>-3194 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1259,-3194,-1258,-3194</points>
<connection>
<GID>2312</GID>
<name>OUT</name></connection>
<intersection>-1258 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1258,-3200.5,-1256.5,-3200.5</points>
<connection>
<GID>2284</GID>
<name>J</name></connection>
<intersection>-1258 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1258,-3204.5,-1256.5,-3204.5</points>
<connection>
<GID>2284</GID>
<name>K</name></connection>
<intersection>-1258 0</intersection></hsegment></shape></wire>
<wire>
<ID>2507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1329,-3199.5,-1321.5,-3199.5</points>
<connection>
<GID>2276</GID>
<name>Q</name></connection>
<connection>
<GID>2277</GID>
<name>J</name></connection>
<intersection>-1328 3</intersection>
<intersection>-1325.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1328,-3234.5,-1328,-3199.5</points>
<intersection>-3234.5 10</intersection>
<intersection>-3219 4</intersection>
<intersection>-3203.5 9</intersection>
<intersection>-3199.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1328,-3219,-1241,-3219</points>
<connection>
<GID>2291</GID>
<name>IN_0</name></connection>
<intersection>-1328 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-1325.5,-3199.5,-1325.5,-3190</points>
<intersection>-3199.5 1</intersection>
<intersection>-3190 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1325.5,-3190,-1314.5,-3190</points>
<connection>
<GID>2302</GID>
<name>IN_0</name></connection>
<intersection>-1325.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1328,-3203.5,-1321.5,-3203.5</points>
<connection>
<GID>2277</GID>
<name>K</name></connection>
<intersection>-1328 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-1328,-3234.5,-1326,-3234.5</points>
<connection>
<GID>2321</GID>
<name>IN_0</name></connection>
<intersection>-1328 3</intersection></hsegment></shape></wire>
<wire>
<ID>2508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1341,-3209,-1075.5,-3209</points>
<intersection>-1341 3</intersection>
<intersection>-1325.5 4</intersection>
<intersection>-1309.5 32</intersection>
<intersection>-1308.5 5</intersection>
<intersection>-1295 31</intersection>
<intersection>-1292.5 16</intersection>
<intersection>-1278 30</intersection>
<intersection>-1276 15</intersection>
<intersection>-1262 29</intersection>
<intersection>-1261 18</intersection>
<intersection>-1244 28</intersection>
<intersection>-1075.5 35</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1341,-3237.5,-1341,-3201.5</points>
<intersection>-3237.5 33</intersection>
<intersection>-3214 39</intersection>
<intersection>-3209 1</intersection>
<intersection>-3201.5 13</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1325.5,-3209,-1325.5,-3201.5</points>
<intersection>-3209 1</intersection>
<intersection>-3201.5 14</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-1308.5,-3209,-1308.5,-3201.5</points>
<intersection>-3209 1</intersection>
<intersection>-3201.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1308.5,-3201.5,-1305.5,-3201.5</points>
<connection>
<GID>2279</GID>
<name>clock</name></connection>
<intersection>-1308.5 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-1341,-3201.5,-1335,-3201.5</points>
<connection>
<GID>2276</GID>
<name>clock</name></connection>
<intersection>-1341 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-1325.5,-3201.5,-1321.5,-3201.5</points>
<connection>
<GID>2277</GID>
<name>clock</name></connection>
<intersection>-1325.5 4</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-1276,-3209,-1276,-3202.5</points>
<intersection>-3209 1</intersection>
<intersection>-3202.5 21</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-1292.5,-3209,-1292.5,-3202</points>
<intersection>-3209 1</intersection>
<intersection>-3202 19</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-1261,-3209,-1261,-3202.5</points>
<intersection>-3209 1</intersection>
<intersection>-3202.5 20</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-1292.5,-3202,-1289.5,-3202</points>
<connection>
<GID>2281</GID>
<name>clock</name></connection>
<intersection>-1292.5 16</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-1261,-3202.5,-1256.5,-3202.5</points>
<connection>
<GID>2284</GID>
<name>clock</name></connection>
<intersection>-1261 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-1276,-3202.5,-1273.5,-3202.5</points>
<connection>
<GID>2283</GID>
<name>clock</name></connection>
<intersection>-1276 15</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-1244,-3237.5,-1244,-3209</points>
<connection>
<GID>2326</GID>
<name>clock</name></connection>
<intersection>-3209 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>-1262,-3237.5,-1262,-3209</points>
<connection>
<GID>2325</GID>
<name>clock</name></connection>
<intersection>-3209 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-1278,-3237.5,-1278,-3209</points>
<connection>
<GID>2324</GID>
<name>clock</name></connection>
<intersection>-3209 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-1295,-3237.5,-1295,-3209</points>
<connection>
<GID>2323</GID>
<name>clock</name></connection>
<intersection>-3209 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-1309.5,-3237.5,-1309.5,-3209</points>
<connection>
<GID>2322</GID>
<name>clock</name></connection>
<intersection>-3209 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-1341,-3237.5,-1326,-3237.5</points>
<connection>
<GID>2321</GID>
<name>clock</name></connection>
<intersection>-1341 3</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>-1075.5,-3276.5,-1075.5,-3209</points>
<intersection>-3276.5 36</intersection>
<intersection>-3209 1</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>-1088.5,-3276.5,-1075.5,-3276.5</points>
<connection>
<GID>2257</GID>
<name>clock</name></connection>
<intersection>-1075.5 35</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-1341.5,-3214,-1341,-3214</points>
<connection>
<GID>2270</GID>
<name>OUT</name></connection>
<intersection>-1341 3</intersection></hsegment></shape></wire>
<wire>
<ID>2509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1314.5,-3234.5,-1314.5,-3192</points>
<connection>
<GID>2302</GID>
<name>IN_1</name></connection>
<intersection>-3234.5 8</intersection>
<intersection>-3218 1</intersection>
<intersection>-3199.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1314.5,-3218,-1241,-3218</points>
<connection>
<GID>2291</GID>
<name>IN_1</name></connection>
<intersection>-1314.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-1315.5,-3199.5,-1314.5,-3199.5</points>
<connection>
<GID>2277</GID>
<name>Q</name></connection>
<intersection>-1314.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1314.5,-3234.5,-1309.5,-3234.5</points>
<connection>
<GID>2322</GID>
<name>IN_0</name></connection>
<intersection>-1314.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1282.5,-3216,-1241,-3216</points>
<connection>
<GID>2291</GID>
<name>IN_3</name></connection>
<intersection>-1282.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1282.5,-3234.5,-1282.5,-3190</points>
<connection>
<GID>2309</GID>
<name>IN_1</name></connection>
<intersection>-3234.5 9</intersection>
<intersection>-3216 1</intersection>
<intersection>-3200 4</intersection>
<intersection>-3190 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1283.5,-3200,-1282.5,-3200</points>
<connection>
<GID>2281</GID>
<name>Q</name></connection>
<intersection>-1282.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1282.5,-3190,-1243,-3190</points>
<connection>
<GID>2315</GID>
<name>IN_1</name></connection>
<intersection>-1282.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1282.5,-3234.5,-1278,-3234.5</points>
<connection>
<GID>2324</GID>
<name>IN_0</name></connection>
<intersection>-1282.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1298.5,-3234.5,-1298.5,-3188</points>
<intersection>-3234.5 9</intersection>
<intersection>-3217 4</intersection>
<intersection>-3199.5 3</intersection>
<intersection>-3193 2</intersection>
<intersection>-3188 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1298.5,-3193,-1297.5,-3193</points>
<connection>
<GID>2306</GID>
<name>IN_1</name></connection>
<intersection>-1298.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1299.5,-3199.5,-1298.5,-3199.5</points>
<connection>
<GID>2279</GID>
<name>Q</name></connection>
<intersection>-1298.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1298.5,-3217,-1241,-3217</points>
<connection>
<GID>2291</GID>
<name>IN_2</name></connection>
<intersection>-1298.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1298.5,-3188,-1243,-3188</points>
<connection>
<GID>2315</GID>
<name>IN_0</name></connection>
<intersection>-1298.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1298.5,-3234.5,-1295,-3234.5</points>
<connection>
<GID>2323</GID>
<name>IN_0</name></connection>
<intersection>-1298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1266.5,-3234.5,-1266.5,-3192</points>
<intersection>-3234.5 8</intersection>
<intersection>-3215 3</intersection>
<intersection>-3200.5 1</intersection>
<intersection>-3192 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1267.5,-3200.5,-1266.5,-3200.5</points>
<connection>
<GID>2283</GID>
<name>Q</name></connection>
<intersection>-1266.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1266.5,-3192,-1243,-3192</points>
<connection>
<GID>2315</GID>
<name>IN_2</name></connection>
<intersection>-1266.5 0</intersection>
<intersection>-1265 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1266.5,-3215,-1241,-3215</points>
<connection>
<GID>2291</GID>
<name>IN_4</name></connection>
<intersection>-1266.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1265,-3195,-1265,-3192</points>
<connection>
<GID>2312</GID>
<name>IN_1</name></connection>
<intersection>-3192 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1266.5,-3234.5,-1262,-3234.5</points>
<connection>
<GID>2325</GID>
<name>IN_0</name></connection>
<intersection>-1266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1248.5,-3234.5,-1248.5,-3194</points>
<intersection>-3234.5 5</intersection>
<intersection>-3214 2</intersection>
<intersection>-3200.5 1</intersection>
<intersection>-3194 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1250.5,-3200.5,-1248.5,-3200.5</points>
<connection>
<GID>2284</GID>
<name>Q</name></connection>
<intersection>-1248.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1248.5,-3214,-1241,-3214</points>
<connection>
<GID>2291</GID>
<name>IN_5</name></connection>
<intersection>-1248.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1248.5,-3194,-1243,-3194</points>
<connection>
<GID>2315</GID>
<name>IN_3</name></connection>
<intersection>-1248.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1248.5,-3234.5,-1244,-3234.5</points>
<connection>
<GID>2326</GID>
<name>IN_0</name></connection>
<intersection>-1248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1318.5,-3249,-1226,-3249</points>
<connection>
<GID>2327</GID>
<name>IN_0</name></connection>
<intersection>-1318.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1318.5,-3258.5,-1318.5,-3234.5</points>
<intersection>-3258.5 8</intersection>
<intersection>-3249 1</intersection>
<intersection>-3234.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1320,-3234.5,-1318.5,-3234.5</points>
<connection>
<GID>2321</GID>
<name>OUT_0</name></connection>
<intersection>-1318.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1320,-3258.5,-1318.5,-3258.5</points>
<connection>
<GID>2274</GID>
<name>IN_3</name></connection>
<intersection>-1318.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2515</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1302,-3248,-1226,-3248</points>
<connection>
<GID>2327</GID>
<name>IN_1</name></connection>
<intersection>-1302 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1302,-3260.5,-1302,-3234.5</points>
<intersection>-3260.5 8</intersection>
<intersection>-3248 1</intersection>
<intersection>-3234.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1303.5,-3234.5,-1302,-3234.5</points>
<connection>
<GID>2322</GID>
<name>OUT_0</name></connection>
<intersection>-1302 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1320,-3260.5,-1302,-3260.5</points>
<connection>
<GID>2274</GID>
<name>IN_2</name></connection>
<intersection>-1302 3</intersection></hsegment></shape></wire>
<wire>
<ID>2516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1288,-3247,-1226,-3247</points>
<connection>
<GID>2327</GID>
<name>IN_2</name></connection>
<intersection>-1288 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1288,-3262.5,-1288,-3234.5</points>
<intersection>-3262.5 8</intersection>
<intersection>-3247 1</intersection>
<intersection>-3234.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1289,-3234.5,-1288,-3234.5</points>
<connection>
<GID>2323</GID>
<name>OUT_0</name></connection>
<intersection>-1288 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1320,-3262.5,-1288,-3262.5</points>
<connection>
<GID>2274</GID>
<name>IN_1</name></connection>
<intersection>-1288 3</intersection></hsegment></shape></wire>
<wire>
<ID>2517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1269.5,-3246,-1226,-3246</points>
<connection>
<GID>2327</GID>
<name>IN_3</name></connection>
<intersection>-1269.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1269.5,-3264.5,-1269.5,-3234.5</points>
<intersection>-3264.5 8</intersection>
<intersection>-3246 1</intersection>
<intersection>-3234.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1272,-3234.5,-1269.5,-3234.5</points>
<connection>
<GID>2324</GID>
<name>OUT_0</name></connection>
<intersection>-1269.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1320,-3264.5,-1269.5,-3264.5</points>
<connection>
<GID>2274</GID>
<name>IN_0</name></connection>
<intersection>-1269.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1288,-3245,-1226,-3245</points>
<connection>
<GID>2327</GID>
<name>IN_4</name></connection>
<intersection>-1288 7</intersection>
<intersection>-1255 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1255,-3245,-1255,-3234.5</points>
<intersection>-3245 1</intersection>
<intersection>-3234.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1256,-3234.5,-1255,-3234.5</points>
<connection>
<GID>2325</GID>
<name>OUT_0</name></connection>
<intersection>-1255 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-1288,-3269,-1288,-3245</points>
<connection>
<GID>2272</GID>
<name>IN_1</name></connection>
<intersection>-3245 1</intersection></vsegment></shape></wire>
<wire>
<ID>2519</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1235,-3244,-1226,-3244</points>
<connection>
<GID>2327</GID>
<name>IN_5</name></connection>
<intersection>-1235 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-1235,-3271,-1235,-3234.5</points>
<intersection>-3271 8</intersection>
<intersection>-3244 1</intersection>
<intersection>-3234.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1238,-3234.5,-1235,-3234.5</points>
<connection>
<GID>2326</GID>
<name>OUT_0</name></connection>
<intersection>-1235 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1288,-3271,-1235,-3271</points>
<connection>
<GID>2272</GID>
<name>IN_0</name></connection>
<intersection>-1235 5</intersection></hsegment></shape></wire>
<wire>
<ID>2520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1178.5,-3276.5,-1178.5,-3264</points>
<intersection>-3276.5 4</intersection>
<intersection>-3272.5 2</intersection>
<intersection>-3264 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1180,-3264,-1169,-3264</points>
<connection>
<GID>2304</GID>
<name>OUT</name></connection>
<connection>
<GID>2305</GID>
<name>IN_0</name></connection>
<intersection>-1178.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1178.5,-3272.5,-1177,-3272.5</points>
<connection>
<GID>2292</GID>
<name>J</name></connection>
<intersection>-1178.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1178.5,-3276.5,-1177,-3276.5</points>
<connection>
<GID>2292</GID>
<name>K</name></connection>
<intersection>-1178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1162,-3277,-1162,-3265</points>
<intersection>-3277 4</intersection>
<intersection>-3273 2</intersection>
<intersection>-3265 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1163,-3265,-1154,-3265</points>
<connection>
<GID>2307</GID>
<name>IN_0</name></connection>
<connection>
<GID>2305</GID>
<name>OUT</name></connection>
<intersection>-1162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1162,-3273,-1161,-3273</points>
<connection>
<GID>2295</GID>
<name>J</name></connection>
<intersection>-1162 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1162,-3277,-1161,-3277</points>
<connection>
<GID>2295</GID>
<name>K</name></connection>
<intersection>-1162 0</intersection></hsegment></shape></wire>
<wire>
<ID>2522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1146.5,-3276.5,-1146.5,-3266</points>
<intersection>-3276.5 4</intersection>
<intersection>-3272.5 2</intersection>
<intersection>-3266 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1148,-3266,-1136.5,-3266</points>
<connection>
<GID>2307</GID>
<name>OUT</name></connection>
<connection>
<GID>2308</GID>
<name>IN_0</name></connection>
<intersection>-1146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1146.5,-3272.5,-1145,-3272.5</points>
<connection>
<GID>2298</GID>
<name>J</name></connection>
<intersection>-1146.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1146.5,-3276.5,-1145,-3276.5</points>
<connection>
<GID>2298</GID>
<name>K</name></connection>
<intersection>-1146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1129.5,-3276.5,-1129.5,-3267</points>
<intersection>-3276.5 4</intersection>
<intersection>-3272.5 2</intersection>
<intersection>-3267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1130.5,-3267,-1129.5,-3267</points>
<connection>
<GID>2308</GID>
<name>OUT</name></connection>
<intersection>-1129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1129.5,-3272.5,-1128,-3272.5</points>
<connection>
<GID>2300</GID>
<name>J</name></connection>
<intersection>-1129.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1129.5,-3276.5,-1128,-3276.5</points>
<connection>
<GID>2300</GID>
<name>K</name></connection>
<intersection>-1129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1200.5,-3272.5,-1193,-3272.5</points>
<connection>
<GID>2288</GID>
<name>Q</name></connection>
<connection>
<GID>2290</GID>
<name>J</name></connection>
<intersection>-1199.5 3</intersection>
<intersection>-1197 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1199.5,-3307.5,-1199.5,-3272.5</points>
<intersection>-3307.5 10</intersection>
<intersection>-3292 4</intersection>
<intersection>-3276.5 9</intersection>
<intersection>-3272.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1199.5,-3292,-1118,-3292</points>
<connection>
<GID>2301</GID>
<name>IN_0</name></connection>
<intersection>-1199.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-1197,-3272.5,-1197,-3263</points>
<intersection>-3272.5 1</intersection>
<intersection>-3263 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1197,-3263,-1186,-3263</points>
<connection>
<GID>2304</GID>
<name>IN_0</name></connection>
<intersection>-1197 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1199.5,-3276.5,-1193,-3276.5</points>
<connection>
<GID>2290</GID>
<name>K</name></connection>
<intersection>-1199.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-1199.5,-3307.5,-1197.5,-3307.5</points>
<connection>
<GID>2311</GID>
<name>IN_0</name></connection>
<intersection>-1199.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1186,-3307.5,-1186,-3265</points>
<connection>
<GID>2304</GID>
<name>IN_1</name></connection>
<intersection>-3307.5 8</intersection>
<intersection>-3291 1</intersection>
<intersection>-3272.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1186,-3291,-1118,-3291</points>
<connection>
<GID>2301</GID>
<name>IN_1</name></connection>
<intersection>-1186 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-1187,-3272.5,-1186,-3272.5</points>
<connection>
<GID>2290</GID>
<name>Q</name></connection>
<intersection>-1186 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1186,-3307.5,-1181,-3307.5</points>
<connection>
<GID>2313</GID>
<name>IN_0</name></connection>
<intersection>-1186 0</intersection></hsegment></shape></wire>
<wire>
<ID>2526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1154,-3289,-1118,-3289</points>
<connection>
<GID>2301</GID>
<name>IN_3</name></connection>
<intersection>-1154 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1154,-3307.5,-1154,-3263</points>
<connection>
<GID>2307</GID>
<name>IN_1</name></connection>
<intersection>-3307.5 9</intersection>
<intersection>-3289 1</intersection>
<intersection>-3273 4</intersection>
<intersection>-3263 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1155,-3273,-1154,-3273</points>
<connection>
<GID>2295</GID>
<name>Q</name></connection>
<intersection>-1154 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1154,-3263,-1114.5,-3263</points>
<connection>
<GID>2310</GID>
<name>IN_1</name></connection>
<intersection>-1154 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1154,-3307.5,-1149.5,-3307.5</points>
<connection>
<GID>2316</GID>
<name>IN_0</name></connection>
<intersection>-1154 3</intersection></hsegment></shape></wire>
<wire>
<ID>2527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1170,-3307.5,-1170,-3261</points>
<intersection>-3307.5 9</intersection>
<intersection>-3290 4</intersection>
<intersection>-3272.5 3</intersection>
<intersection>-3266 2</intersection>
<intersection>-3261 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1170,-3266,-1169,-3266</points>
<connection>
<GID>2305</GID>
<name>IN_1</name></connection>
<intersection>-1170 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1171,-3272.5,-1170,-3272.5</points>
<connection>
<GID>2292</GID>
<name>Q</name></connection>
<intersection>-1170 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-1170,-3290,-1118,-3290</points>
<connection>
<GID>2301</GID>
<name>IN_2</name></connection>
<intersection>-1170 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-1170,-3261,-1114.5,-3261</points>
<connection>
<GID>2310</GID>
<name>IN_0</name></connection>
<intersection>-1170 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1170,-3307.5,-1166.5,-3307.5</points>
<connection>
<GID>2314</GID>
<name>IN_0</name></connection>
<intersection>-1170 0</intersection></hsegment></shape></wire>
<wire>
<ID>2528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1138,-3307.5,-1138,-3265</points>
<intersection>-3307.5 8</intersection>
<intersection>-3288 3</intersection>
<intersection>-3272.5 1</intersection>
<intersection>-3265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1139,-3272.5,-1138,-3272.5</points>
<connection>
<GID>2298</GID>
<name>Q</name></connection>
<intersection>-1138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1138,-3265,-1114.5,-3265</points>
<connection>
<GID>2310</GID>
<name>IN_2</name></connection>
<intersection>-1138 0</intersection>
<intersection>-1136.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1138,-3288,-1118,-3288</points>
<connection>
<GID>2301</GID>
<name>IN_4</name></connection>
<intersection>-1138 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1136.5,-3268,-1136.5,-3265</points>
<connection>
<GID>2308</GID>
<name>IN_1</name></connection>
<intersection>-3265 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1138,-3307.5,-1133.5,-3307.5</points>
<connection>
<GID>2317</GID>
<name>IN_0</name></connection>
<intersection>-1138 0</intersection></hsegment></shape></wire>
<wire>
<ID>2529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1120,-3307.5,-1120,-3267</points>
<intersection>-3307.5 5</intersection>
<intersection>-3287 2</intersection>
<intersection>-3272.5 1</intersection>
<intersection>-3267 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1122,-3272.5,-1120,-3272.5</points>
<connection>
<GID>2300</GID>
<name>Q</name></connection>
<intersection>-1120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1120,-3287,-1118,-3287</points>
<connection>
<GID>2301</GID>
<name>IN_5</name></connection>
<intersection>-1120 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-1120,-3267,-1114.5,-3267</points>
<connection>
<GID>2310</GID>
<name>IN_3</name></connection>
<intersection>-1120 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1120,-3307.5,-1115.5,-3307.5</points>
<connection>
<GID>2318</GID>
<name>IN_0</name></connection>
<intersection>-1120 0</intersection></hsegment></shape></wire>
<wire>
<ID>2530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1190,-3359.5,-689,-3359.5</points>
<intersection>-1190 3</intersection>
<intersection>-689 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1190,-3359.5,-1190,-3307.5</points>
<intersection>-3359.5 1</intersection>
<intersection>-3322 7</intersection>
<intersection>-3307.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1191.5,-3307.5,-1190,-3307.5</points>
<connection>
<GID>2311</GID>
<name>OUT_0</name></connection>
<intersection>-1190 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-689,-4930,-689,-3359.5</points>
<intersection>-4930 56</intersection>
<intersection>-4708.5 54</intersection>
<intersection>-4469 53</intersection>
<intersection>-4210.5 52</intersection>
<intersection>-4044 51</intersection>
<intersection>-3862 50</intersection>
<intersection>-3713 49</intersection>
<intersection>-3586 23</intersection>
<intersection>-3359.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1190,-3322,-1097.5,-3322</points>
<connection>
<GID>2319</GID>
<name>IN_0</name></connection>
<intersection>-1190 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-869,-3586,-689,-3586</points>
<intersection>-869 29</intersection>
<intersection>-689 5</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>-869,-3589.5,-869,-3586</points>
<connection>
<GID>2331</GID>
<name>IN_0</name></connection>
<intersection>-3586 23</intersection></vsegment>
<hsegment>
<ID>49</ID>
<points>-779,-3713,-689,-3713</points>
<connection>
<GID>2376</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-777.5,-3862,-689,-3862</points>
<connection>
<GID>1873</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>-775,-4044,-689,-4044</points>
<connection>
<GID>1939</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>-762.5,-4210.5,-689,-4210.5</points>
<connection>
<GID>1973</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>-771.5,-4469,-689,-4469</points>
<connection>
<GID>1991</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>-771,-4708.5,-689,-4708.5</points>
<connection>
<GID>2036</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>-753.5,-4930,-689,-4930</points>
<connection>
<GID>2059</GID>
<name>IN_0</name></connection>
<intersection>-689 5</intersection></hsegment></shape></wire>
<wire>
<ID>2531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1173.5,-3355,-692.5,-3355</points>
<intersection>-1173.5 3</intersection>
<intersection>-692.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1173.5,-3355,-1173.5,-3307.5</points>
<intersection>-3355 1</intersection>
<intersection>-3321 7</intersection>
<intersection>-3307.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1175,-3307.5,-1173.5,-3307.5</points>
<connection>
<GID>2313</GID>
<name>OUT_0</name></connection>
<intersection>-1173.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-692.5,-4921.5,-692.5,-3355</points>
<intersection>-4921.5 56</intersection>
<intersection>-4699 54</intersection>
<intersection>-4463 53</intersection>
<intersection>-4202 30</intersection>
<intersection>-4032 52</intersection>
<intersection>-3856.5 51</intersection>
<intersection>-3710 50</intersection>
<intersection>-3584 19</intersection>
<intersection>-3355 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1173.5,-3321,-1097.5,-3321</points>
<connection>
<GID>2319</GID>
<name>IN_1</name></connection>
<intersection>-1173.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-855.5,-3584,-692.5,-3584</points>
<intersection>-855.5 25</intersection>
<intersection>-692.5 5</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-855.5,-3589.5,-855.5,-3584</points>
<connection>
<GID>2332</GID>
<name>IN_0</name></connection>
<intersection>-3584 19</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>-750.5,-4202,-692.5,-4202</points>
<connection>
<GID>1975</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-765.5,-3710,-692.5,-3710</points>
<connection>
<GID>2378</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>-762,-3856.5,-692.5,-3856.5</points>
<connection>
<GID>1877</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>-765,-4032,-692.5,-4032</points>
<connection>
<GID>1958</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>-760.5,-4463,-692.5,-4463</points>
<connection>
<GID>1992</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>-760,-4699,-692.5,-4699</points>
<connection>
<GID>2038</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>-741.5,-4921.5,-692.5,-4921.5</points>
<connection>
<GID>2062</GID>
<name>IN_0</name></connection>
<intersection>-692.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>2532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1159.5,-3350.5,-695,-3350.5</points>
<intersection>-1159.5 3</intersection>
<intersection>-695 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1159.5,-3350.5,-1159.5,-3307.5</points>
<intersection>-3350.5 1</intersection>
<intersection>-3320 7</intersection>
<intersection>-3307.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1160.5,-3307.5,-1159.5,-3307.5</points>
<connection>
<GID>2314</GID>
<name>OUT_0</name></connection>
<intersection>-1159.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-695,-4911.5,-695,-3350.5</points>
<intersection>-4911.5 52</intersection>
<intersection>-4689.5 50</intersection>
<intersection>-4453.5 49</intersection>
<intersection>-4192 48</intersection>
<intersection>-4023.5 47</intersection>
<intersection>-3848.5 21</intersection>
<intersection>-3702.5 46</intersection>
<intersection>-3581.5 19</intersection>
<intersection>-3350.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1159.5,-3320,-1097.5,-3320</points>
<connection>
<GID>2319</GID>
<name>IN_2</name></connection>
<intersection>-1159.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-842.5,-3581.5,-695,-3581.5</points>
<intersection>-842.5 25</intersection>
<intersection>-695 5</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-761.5,-3848.5,-695,-3848.5</points>
<connection>
<GID>1882</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-842.5,-3589.5,-842.5,-3581.5</points>
<connection>
<GID>2334</GID>
<name>IN_0</name></connection>
<intersection>-3581.5 19</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>-766,-3702.5,-695,-3702.5</points>
<connection>
<GID>2381</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>-765,-4023.5,-695,-4023.5</points>
<connection>
<GID>1959</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-750.5,-4192,-695,-4192</points>
<connection>
<GID>1976</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>-760.5,-4453.5,-695,-4453.5</points>
<connection>
<GID>2013</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-760.5,-4689.5,-695,-4689.5</points>
<connection>
<GID>2040</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>-740,-4911.5,-695,-4911.5</points>
<connection>
<GID>2064</GID>
<name>IN_0</name></connection>
<intersection>-695 5</intersection></hsegment></shape></wire>
<wire>
<ID>2533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1141,-3346,-697,-3346</points>
<intersection>-1141 3</intersection>
<intersection>-697 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1141,-3346,-1141,-3307.5</points>
<intersection>-3346 1</intersection>
<intersection>-3319 7</intersection>
<intersection>-3307.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1143.5,-3307.5,-1141,-3307.5</points>
<connection>
<GID>2316</GID>
<name>OUT_0</name></connection>
<intersection>-1141 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-697,-4902,-697,-3346</points>
<intersection>-4902 53</intersection>
<intersection>-4681 51</intersection>
<intersection>-4444 50</intersection>
<intersection>-4185 49</intersection>
<intersection>-4016 48</intersection>
<intersection>-3840.5 23</intersection>
<intersection>-3694.5 47</intersection>
<intersection>-3579 21</intersection>
<intersection>-3346 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1141,-3319,-1097.5,-3319</points>
<connection>
<GID>2319</GID>
<name>IN_3</name></connection>
<intersection>-1141 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-829.5,-3579,-697,-3579</points>
<intersection>-829.5 27</intersection>
<intersection>-697 5</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-760.5,-3840.5,-697,-3840.5</points>
<connection>
<GID>1887</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>-829.5,-3589.5,-829.5,-3579</points>
<connection>
<GID>2336</GID>
<name>IN_0</name></connection>
<intersection>-3579 21</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>-765,-3694.5,-697,-3694.5</points>
<connection>
<GID>2383</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-764,-4016,-697,-4016</points>
<connection>
<GID>1962</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>-749,-4185,-697,-4185</points>
<connection>
<GID>1978</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-759.5,-4444,-697,-4444</points>
<connection>
<GID>2016</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>-760,-4681,-697,-4681</points>
<connection>
<GID>2042</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>-739.5,-4902,-697,-4902</points>
<connection>
<GID>2118</GID>
<name>IN_0</name></connection>
<intersection>-697 5</intersection></hsegment></shape></wire>
<wire>
<ID>2534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1126,-3343,-701,-3343</points>
<intersection>-1126 3</intersection>
<intersection>-701 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1126,-3343,-1126,-3307.5</points>
<intersection>-3343 1</intersection>
<intersection>-3318 7</intersection>
<intersection>-3307.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1127.5,-3307.5,-1126,-3307.5</points>
<connection>
<GID>2317</GID>
<name>OUT_0</name></connection>
<intersection>-1126 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-701,-4893.5,-701,-3343</points>
<intersection>-4893.5 49</intersection>
<intersection>-4672.5 47</intersection>
<intersection>-4435.5 46</intersection>
<intersection>-4175.5 45</intersection>
<intersection>-4007 44</intersection>
<intersection>-3830 19</intersection>
<intersection>-3688.5 43</intersection>
<intersection>-3576 17</intersection>
<intersection>-3343 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1126,-3318,-1097.5,-3318</points>
<connection>
<GID>2319</GID>
<name>IN_4</name></connection>
<intersection>-1126 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-817,-3576,-701,-3576</points>
<intersection>-817 23</intersection>
<intersection>-701 5</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-760,-3830,-701,-3830</points>
<connection>
<GID>1889</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-817,-3590,-817,-3576</points>
<connection>
<GID>2337</GID>
<name>IN_0</name></connection>
<intersection>-3576 17</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>-765,-3688.5,-701,-3688.5</points>
<connection>
<GID>2385</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>-763.5,-4007,-701,-4007</points>
<connection>
<GID>1964</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-748.5,-4175.5,-701,-4175.5</points>
<connection>
<GID>1980</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>-759,-4435.5,-701,-4435.5</points>
<connection>
<GID>2029</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>-760,-4672.5,-701,-4672.5</points>
<connection>
<GID>2044</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>-740,-4893.5,-701,-4893.5</points>
<connection>
<GID>2125</GID>
<name>IN_0</name></connection>
<intersection>-701 5</intersection></hsegment></shape></wire>
<wire>
<ID>2535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1103.5,-3338,-1103.5,-3307.5</points>
<intersection>-3338 5</intersection>
<intersection>-3317 8</intersection>
<intersection>-3307.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1109.5,-3307.5,-1103.5,-3307.5</points>
<connection>
<GID>2318</GID>
<name>OUT_0</name></connection>
<intersection>-1103.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-1103.5,-3338,-705.5,-3338</points>
<intersection>-1103.5 0</intersection>
<intersection>-705.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-705.5,-4885,-705.5,-3338</points>
<intersection>-4885 50</intersection>
<intersection>-4665 48</intersection>
<intersection>-4427 47</intersection>
<intersection>-4168.5 46</intersection>
<intersection>-3999 45</intersection>
<intersection>-3819 20</intersection>
<intersection>-3683 44</intersection>
<intersection>-3572 18</intersection>
<intersection>-3338 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1103.5,-3317,-1097.5,-3317</points>
<connection>
<GID>2319</GID>
<name>IN_5</name></connection>
<intersection>-1103.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-804.5,-3572,-705.5,-3572</points>
<intersection>-804.5 24</intersection>
<intersection>-705.5 6</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-760.5,-3819,-705.5,-3819</points>
<connection>
<GID>1894</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-804.5,-3590,-804.5,-3572</points>
<connection>
<GID>2339</GID>
<name>IN_0</name></connection>
<intersection>-3572 18</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>-764.5,-3683,-705.5,-3683</points>
<connection>
<GID>2388</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-763,-3999,-705.5,-3999</points>
<connection>
<GID>1966</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>-748,-4168.5,-705.5,-4168.5</points>
<connection>
<GID>1982</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>-758,-4427,-705.5,-4427</points>
<connection>
<GID>2030</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-759.5,-4665,-705.5,-4665</points>
<connection>
<GID>2046</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-740.5,-4885,-705.5,-4885</points>
<connection>
<GID>2303</GID>
<name>IN_0</name></connection>
<intersection>-705.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>2536</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-1210,-3272.5,-1210,-3251.5</points>
<intersection>-3272.5 17</intersection>
<intersection>-3251.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1349,-3251.5,-1088.5,-3251.5</points>
<intersection>-1349 11</intersection>
<intersection>-1210 3</intersection>
<intersection>-1206.5 44</intersection>
<intersection>-1088.5 43</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-1349,-3199.5,-1335,-3199.5</points>
<connection>
<GID>2276</GID>
<name>J</name></connection>
<intersection>-1349 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-1349,-3265,-1349,-3199.5</points>
<intersection>-3265 22</intersection>
<intersection>-3252 23</intersection>
<intersection>-3251.5 4</intersection>
<intersection>-3213 21</intersection>
<intersection>-3205.5 28</intersection>
<intersection>-3203.5 14</intersection>
<intersection>-3199.5 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-1349,-3203.5,-1335,-3203.5</points>
<connection>
<GID>2276</GID>
<name>K</name></connection>
<intersection>-1349 11</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-1210,-3272.5,-1206.5,-3272.5</points>
<connection>
<GID>2288</GID>
<name>J</name></connection>
<intersection>-1210 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-1349,-3213,-1347.5,-3213</points>
<connection>
<GID>2270</GID>
<name>IN_0</name></connection>
<intersection>-1349 11</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-1351.5,-3265,-1349,-3265</points>
<connection>
<GID>2289</GID>
<name>IN_1</name></connection>
<intersection>-1349 11</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-1349,-3252,-1340.5,-3252</points>
<intersection>-1349 11</intersection>
<intersection>-1340.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-1340.5,-3256.5,-1340.5,-3252</points>
<connection>
<GID>2278</GID>
<name>IN_1</name></connection>
<intersection>-3252 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-1355.5,-3205.5,-1349,-3205.5</points>
<connection>
<GID>2328</GID>
<name>OUT</name></connection>
<intersection>-1349 11</intersection></hsegment>
<vsegment>
<ID>43</ID>
<points>-1088.5,-3278.5,-1088.5,-3251.5</points>
<connection>
<GID>2257</GID>
<name>J</name></connection>
<intersection>-3251.5 4</intersection></vsegment>
<vsegment>
<ID>44</ID>
<points>-1206.5,-3276.5,-1206.5,-3251.5</points>
<connection>
<GID>2288</GID>
<name>K</name></connection>
<intersection>-3251.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>2537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1207.5,-3310.5,-1207.5,-3219.5</points>
<intersection>-3310.5 8</intersection>
<intersection>-3274.5 1</intersection>
<intersection>-3219.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1207.5,-3274.5,-1128,-3274.5</points>
<connection>
<GID>2288</GID>
<name>clock</name></connection>
<connection>
<GID>2290</GID>
<name>clock</name></connection>
<connection>
<GID>2292</GID>
<name>clock</name></connection>
<connection>
<GID>2298</GID>
<name>clock</name></connection>
<connection>
<GID>2300</GID>
<name>clock</name></connection>
<intersection>-1207.5 0</intersection>
<intersection>-1161 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1161,-3275,-1161,-3274.5</points>
<connection>
<GID>2295</GID>
<name>clock</name></connection>
<intersection>-3274.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1207.5,-3310.5,-1115.5,-3310.5</points>
<connection>
<GID>2311</GID>
<name>clock</name></connection>
<connection>
<GID>2313</GID>
<name>clock</name></connection>
<connection>
<GID>2314</GID>
<name>clock</name></connection>
<connection>
<GID>2316</GID>
<name>clock</name></connection>
<connection>
<GID>2317</GID>
<name>clock</name></connection>
<connection>
<GID>2318</GID>
<name>clock</name></connection>
<intersection>-1207.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-1207.5,-3219.5,-1205,-3219.5</points>
<connection>
<GID>2320</GID>
<name>OUT_0</name></connection>
<intersection>-1207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-822.5,-4506,-822.5,-4501</points>
<connection>
<GID>2172</GID>
<name>OUT_0</name></connection>
<intersection>-4506 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-820.5,-4512.5,-820.5,-4506</points>
<connection>
<GID>2246</GID>
<name>IN_2</name></connection>
<intersection>-4506 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-822.5,-4506,-820.5,-4506</points>
<intersection>-822.5 0</intersection>
<intersection>-820.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-807.5,-4506.5,-807.5,-4501</points>
<connection>
<GID>2173</GID>
<name>OUT_0</name></connection>
<intersection>-4506.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-818.5,-4512.5,-818.5,-4506.5</points>
<connection>
<GID>2246</GID>
<name>IN_1</name></connection>
<intersection>-4506.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-818.5,-4506.5,-807.5,-4506.5</points>
<intersection>-818.5 1</intersection>
<intersection>-807.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-796,-4507.5,-796,-4500.5</points>
<connection>
<GID>2176</GID>
<name>OUT_0</name></connection>
<intersection>-4507.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-816.5,-4512.5,-816.5,-4507.5</points>
<connection>
<GID>2246</GID>
<name>IN_0</name></connection>
<intersection>-4507.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-816.5,-4507.5,-796,-4507.5</points>
<intersection>-816.5 1</intersection>
<intersection>-796 0</intersection></hsegment></shape></wire>
<wire>
<ID>2541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-783,-4506,-783,-4501</points>
<connection>
<GID>2178</GID>
<name>OUT_0</name></connection>
<intersection>-4506 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-784,-4511.5,-784,-4506</points>
<connection>
<GID>2343</GID>
<name>IN_1</name></connection>
<intersection>-4506 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-784,-4506,-783,-4506</points>
<intersection>-784 1</intersection>
<intersection>-783 0</intersection></hsegment></shape></wire>
<wire>
<ID>2542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-770,-4506,-770,-4500.5</points>
<connection>
<GID>2179</GID>
<name>OUT_0</name></connection>
<intersection>-4506 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-782,-4511.5,-782,-4506</points>
<connection>
<GID>2343</GID>
<name>IN_0</name></connection>
<intersection>-4506 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-782,-4506,-770,-4506</points>
<intersection>-782 1</intersection>
<intersection>-770 0</intersection></hsegment></shape></wire>
<wire>
<ID>2543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-819.5,-4522,-819.5,-4518.5</points>
<connection>
<GID>2246</GID>
<name>OUT</name></connection>
<intersection>-4522 8</intersection>
<intersection>-4521.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-806.5,-4534.5,-806.5,-4521.5</points>
<connection>
<GID>2345</GID>
<name>IN_1</name></connection>
<intersection>-4529.5 7</intersection>
<intersection>-4521.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-819.5,-4521.5,-806.5,-4521.5</points>
<intersection>-819.5 0</intersection>
<intersection>-806.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-806.5,-4529.5,-795,-4529.5</points>
<connection>
<GID>2382</GID>
<name>IN_0</name></connection>
<intersection>-806.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-870,-4522,-819.5,-4522</points>
<connection>
<GID>1960</GID>
<name>IN_0</name></connection>
<intersection>-819.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-985,-3769.5,-985,-3655</points>
<connection>
<GID>2074</GID>
<name>OUT</name></connection>
<intersection>-3769.5 13</intersection>
<intersection>-3709 1</intersection>
<intersection>-3700.5 7</intersection>
<intersection>-3692 3</intersection>
<intersection>-3684 8</intersection>
<intersection>-3675.5 5</intersection>
<intersection>-3662.5 15</intersection>
<intersection>-3657.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-985,-3709,-962,-3709</points>
<connection>
<GID>2346</GID>
<name>IN_0</name></connection>
<intersection>-985 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-985,-3692,-963,-3692</points>
<connection>
<GID>2348</GID>
<name>IN_0</name></connection>
<intersection>-985 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-985,-3675.5,-964,-3675.5</points>
<connection>
<GID>2350</GID>
<name>IN_0</name></connection>
<intersection>-985 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-985,-3700.5,-962.5,-3700.5</points>
<connection>
<GID>2347</GID>
<name>IN_0</name></connection>
<intersection>-985 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-985,-3684,-963.5,-3684</points>
<connection>
<GID>2349</GID>
<name>IN_0</name></connection>
<intersection>-985 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-985,-3657.5,-964,-3657.5</points>
<intersection>-985 0</intersection>
<intersection>-964 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-964,-3667,-964,-3657.5</points>
<connection>
<GID>2351</GID>
<name>IN_0</name></connection>
<intersection>-3657.5 9</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-985,-3769.5,-774.5,-3769.5</points>
<intersection>-985 0</intersection>
<intersection>-774.5 16</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-985,-3662.5,-784,-3662.5</points>
<connection>
<GID>2373</GID>
<name>IN_1</name></connection>
<intersection>-985 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-774.5,-3769.5,-774.5,-3765</points>
<connection>
<GID>1867</GID>
<name>IN_1</name></connection>
<intersection>-3769.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>2545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-783,-4521,-783,-4517.5</points>
<connection>
<GID>2343</GID>
<name>OUT</name></connection>
<intersection>-4521 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-804.5,-4534.5,-804.5,-4521</points>
<connection>
<GID>2345</GID>
<name>IN_0</name></connection>
<intersection>-4531.5 6</intersection>
<intersection>-4524 7</intersection>
<intersection>-4521 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-804.5,-4521,-783,-4521</points>
<intersection>-804.5 1</intersection>
<intersection>-783 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-804.5,-4531.5,-795,-4531.5</points>
<connection>
<GID>2382</GID>
<name>IN_1</name></connection>
<intersection>-804.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-910.5,-4524,-804.5,-4524</points>
<connection>
<GID>1906</GID>
<name>IN_0</name></connection>
<intersection>-804.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-931.5,-4443.5,-872.5,-4443.5</points>
<connection>
<GID>2394</GID>
<name>OUT</name></connection>
<connection>
<GID>2377</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-849.5,-4479.5,-849.5,-4443.5</points>
<connection>
<GID>2352</GID>
<name>IN_1</name></connection>
<intersection>-4443.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-866.5,-4443.5,-849.5,-4443.5</points>
<connection>
<GID>2377</GID>
<name>Q</name></connection>
<intersection>-849.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-932,-4433.5,-885.5,-4433.5</points>
<connection>
<GID>2396</GID>
<name>OUT</name></connection>
<connection>
<GID>2379</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-836,-4479.5,-836,-4433.5</points>
<connection>
<GID>2354</GID>
<name>IN_1</name></connection>
<intersection>-4433.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-879.5,-4433.5,-836,-4433.5</points>
<connection>
<GID>2379</GID>
<name>Q</name></connection>
<intersection>-836 0</intersection></hsegment></shape></wire>
<wire>
<ID>2550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-933.5,-4422.5,-898.5,-4422.5</points>
<connection>
<GID>2397</GID>
<name>OUT</name></connection>
<connection>
<GID>2380</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-823,-4479.5,-823,-4422.5</points>
<connection>
<GID>2356</GID>
<name>IN_1</name></connection>
<intersection>-4422.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-892.5,-4422.5,-823,-4422.5</points>
<connection>
<GID>2380</GID>
<name>Q</name></connection>
<intersection>-823 0</intersection></hsegment></shape></wire>
<wire>
<ID>2552</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-953,-3553.5,-894,-3553.5</points>
<connection>
<GID>2171</GID>
<name>OUT</name></connection>
<connection>
<GID>2360</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-871,-3589.5,-871,-3553.5</points>
<connection>
<GID>2331</GID>
<name>IN_1</name></connection>
<intersection>-3553.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-888,-3553.5,-871,-3553.5</points>
<connection>
<GID>2360</GID>
<name>Q</name></connection>
<intersection>-871 0</intersection></hsegment></shape></wire>
<wire>
<ID>2554</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-953.5,-3543.5,-907,-3543.5</points>
<connection>
<GID>2174</GID>
<name>OUT</name></connection>
<connection>
<GID>2363</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-857.5,-3589.5,-857.5,-3543.5</points>
<connection>
<GID>2332</GID>
<name>IN_1</name></connection>
<intersection>-3543.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-901,-3543.5,-857.5,-3543.5</points>
<connection>
<GID>2363</GID>
<name>Q</name></connection>
<intersection>-857.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-955,-3532.5,-920,-3532.5</points>
<connection>
<GID>2175</GID>
<name>OUT</name></connection>
<connection>
<GID>2364</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844.5,-3589.5,-844.5,-3532.5</points>
<connection>
<GID>2334</GID>
<name>IN_1</name></connection>
<intersection>-3532.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-914,-3532.5,-844.5,-3532.5</points>
<connection>
<GID>2364</GID>
<name>Q</name></connection>
<intersection>-844.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2558</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-955.5,-3523.5,-927.5,-3523.5</points>
<connection>
<GID>2177</GID>
<name>OUT</name></connection>
<connection>
<GID>2365</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-831.5,-3589.5,-831.5,-3523.5</points>
<connection>
<GID>2336</GID>
<name>IN_1</name></connection>
<intersection>-3523.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-921.5,-3523.5,-831.5,-3523.5</points>
<connection>
<GID>2365</GID>
<name>Q</name></connection>
<intersection>-831.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2560</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-956.5,-3516,-936,-3516</points>
<connection>
<GID>2180</GID>
<name>OUT</name></connection>
<connection>
<GID>2366</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-819,-3590,-819,-3516</points>
<connection>
<GID>2337</GID>
<name>IN_1</name></connection>
<intersection>-3516 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-930,-3516,-819,-3516</points>
<connection>
<GID>2366</GID>
<name>Q</name></connection>
<intersection>-819 0</intersection></hsegment></shape></wire>
<wire>
<ID>2562</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-957.5,-3508.5,-945,-3508.5</points>
<connection>
<GID>2181</GID>
<name>OUT</name></connection>
<connection>
<GID>2367</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-806.5,-3590,-806.5,-3508.5</points>
<connection>
<GID>2339</GID>
<name>IN_1</name></connection>
<intersection>-3508.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-939,-3508.5,-806.5,-3508.5</points>
<connection>
<GID>2367</GID>
<name>Q</name></connection>
<intersection>-806.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-956,-3710,-904,-3710</points>
<connection>
<GID>2346</GID>
<name>OUT</name></connection>
<connection>
<GID>2368</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-934,-4413.5,-906,-4413.5</points>
<connection>
<GID>2398</GID>
<name>OUT</name></connection>
<connection>
<GID>2384</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-810,-4479.5,-810,-4413.5</points>
<connection>
<GID>2357</GID>
<name>IN_1</name></connection>
<intersection>-4413.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-900,-4413.5,-810,-4413.5</points>
<connection>
<GID>2384</GID>
<name>Q</name></connection>
<intersection>-810 0</intersection></hsegment></shape></wire>
<wire>
<ID>2567</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-935,-4406,-914.5,-4406</points>
<connection>
<GID>2399</GID>
<name>OUT</name></connection>
<connection>
<GID>2386</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-797.5,-4480,-797.5,-4406</points>
<connection>
<GID>2358</GID>
<name>IN_1</name></connection>
<intersection>-4406 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-908.5,-4406,-797.5,-4406</points>
<connection>
<GID>2386</GID>
<name>Q</name></connection>
<intersection>-797.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2569</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-936,-4398.5,-923.5,-4398.5</points>
<connection>
<GID>2400</GID>
<name>OUT</name></connection>
<connection>
<GID>2389</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-785,-4480,-785,-4398.5</points>
<connection>
<GID>2359</GID>
<name>IN_1</name></connection>
<intersection>-4398.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-917.5,-4398.5,-785,-4398.5</points>
<connection>
<GID>2389</GID>
<name>Q</name></connection>
<intersection>-785 0</intersection></hsegment></shape></wire>
<wire>
<ID>2571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-928.5,-4445.5,-928.5,-4394.5</points>
<connection>
<GID>2392</GID>
<name>OUT_0</name></connection>
<intersection>-4445.5 7</intersection>
<intersection>-4435.5 5</intersection>
<intersection>-4424.5 8</intersection>
<intersection>-4415.5 3</intersection>
<intersection>-4408 9</intersection>
<intersection>-4400.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-928.5,-4400.5,-923.5,-4400.5</points>
<connection>
<GID>2389</GID>
<name>clock</name></connection>
<intersection>-928.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-928.5,-4415.5,-906,-4415.5</points>
<connection>
<GID>2384</GID>
<name>clock</name></connection>
<intersection>-928.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-928.5,-4435.5,-885.5,-4435.5</points>
<connection>
<GID>2379</GID>
<name>clock</name></connection>
<intersection>-928.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-928.5,-4445.5,-872.5,-4445.5</points>
<connection>
<GID>2377</GID>
<name>clock</name></connection>
<intersection>-928.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-928.5,-4424.5,-898.5,-4424.5</points>
<connection>
<GID>2380</GID>
<name>clock</name></connection>
<intersection>-928.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-928.5,-4408,-914.5,-4408</points>
<connection>
<GID>2386</GID>
<name>clock</name></connection>
<intersection>-928.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-966.5,-4766.5,-966.5,-4611.5</points>
<connection>
<GID>2122</GID>
<name>OUT</name></connection>
<intersection>-4766.5 13</intersection>
<intersection>-4676.5 1</intersection>
<intersection>-4666.5 3</intersection>
<intersection>-4655.5 5</intersection>
<intersection>-4646.5 7</intersection>
<intersection>-4639 9</intersection>
<intersection>-4615 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-966.5,-4676.5,-935.5,-4676.5</points>
<connection>
<GID>2434</GID>
<name>IN_0</name></connection>
<intersection>-966.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-966.5,-4666.5,-936,-4666.5</points>
<connection>
<GID>2435</GID>
<name>IN_0</name></connection>
<intersection>-966.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-966.5,-4655.5,-937.5,-4655.5</points>
<connection>
<GID>2436</GID>
<name>IN_0</name></connection>
<intersection>-966.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-966.5,-4646.5,-938,-4646.5</points>
<connection>
<GID>2437</GID>
<name>IN_0</name></connection>
<intersection>-966.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-966.5,-4639,-939,-4639</points>
<connection>
<GID>2438</GID>
<name>IN_0</name></connection>
<intersection>-966.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-966.5,-4615,-781,-4615</points>
<intersection>-966.5 0</intersection>
<intersection>-940 15</intersection>
<intersection>-781 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-966.5,-4766.5,-781,-4766.5</points>
<connection>
<GID>1883</GID>
<name>IN_1</name></connection>
<intersection>-966.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-781,-4615,-781,-4552.5</points>
<connection>
<GID>2034</GID>
<name>IN_1</name></connection>
<intersection>-4615 11</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-940,-4631.5,-940,-4615</points>
<connection>
<GID>2439</GID>
<name>IN_0</name></connection>
<intersection>-4615 11</intersection></vsegment></shape></wire>
<wire>
<ID>2573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-846.5,-4723,-846.5,-4719.5</points>
<connection>
<GID>2417</GID>
<name>OUT</name></connection>
<intersection>-4723 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-846.5,-4723,-845.5,-4723</points>
<connection>
<GID>2440</GID>
<name>IN_0</name></connection>
<intersection>-846.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-833,-4723.5,-833,-4719.5</points>
<connection>
<GID>2418</GID>
<name>OUT</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-833,-4723.5,-829.5,-4723.5</points>
<connection>
<GID>2402</GID>
<name>IN_0</name></connection>
<intersection>-833 0</intersection></hsegment></shape></wire>
<wire>
<ID>2575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-820,-4723.5,-820,-4719.5</points>
<connection>
<GID>2419</GID>
<name>OUT</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-820,-4723.5,-816,-4723.5</points>
<connection>
<GID>2403</GID>
<name>IN_0</name></connection>
<intersection>-820 0</intersection></hsegment></shape></wire>
<wire>
<ID>2576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-804,-4723.5,-804,-4719.5</points>
<intersection>-4723.5 1</intersection>
<intersection>-4719.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-804,-4723.5,-801,-4723.5</points>
<connection>
<GID>2404</GID>
<name>IN_0</name></connection>
<intersection>-804 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-807,-4719.5,-804,-4719.5</points>
<connection>
<GID>2420</GID>
<name>OUT</name></connection>
<intersection>-804 0</intersection></hsegment></shape></wire>
<wire>
<ID>2577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-794.5,-4722,-794.5,-4720</points>
<connection>
<GID>2421</GID>
<name>OUT</name></connection>
<intersection>-4722 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-794.5,-4722,-790.5,-4722</points>
<intersection>-794.5 0</intersection>
<intersection>-790.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-790.5,-4723.5,-790.5,-4722</points>
<connection>
<GID>2405</GID>
<name>IN_0</name></connection>
<intersection>-4722 1</intersection></vsegment></shape></wire>
<wire>
<ID>2578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-782,-4722,-782,-4720</points>
<connection>
<GID>2423</GID>
<name>OUT</name></connection>
<intersection>-4722 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-782,-4722,-777.5,-4722</points>
<intersection>-782 0</intersection>
<intersection>-777.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-777.5,-4723.5,-777.5,-4722</points>
<connection>
<GID>2406</GID>
<name>IN_0</name></connection>
<intersection>-4722 1</intersection></vsegment></shape></wire>
<wire>
<ID>2579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-835.5,-4731,-835.5,-4723</points>
<connection>
<GID>2407</GID>
<name>IN_0</name></connection>
<intersection>-4723 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-839.5,-4723,-835.5,-4723</points>
<connection>
<GID>2440</GID>
<name>OUT_0</name></connection>
<intersection>-835.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-820.5,-4731,-820.5,-4723.5</points>
<connection>
<GID>2408</GID>
<name>IN_0</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-823.5,-4723.5,-820.5,-4723.5</points>
<connection>
<GID>2402</GID>
<name>OUT_0</name></connection>
<intersection>-820.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805.5,-4731,-805.5,-4723.5</points>
<connection>
<GID>2409</GID>
<name>IN_0</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-810,-4723.5,-805.5,-4723.5</points>
<connection>
<GID>2403</GID>
<name>OUT_0</name></connection>
<intersection>-805.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2582</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-794,-4730.5,-794,-4723.5</points>
<connection>
<GID>2410</GID>
<name>IN_0</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-795,-4723.5,-794,-4723.5</points>
<connection>
<GID>2404</GID>
<name>OUT_0</name></connection>
<intersection>-794 0</intersection></hsegment></shape></wire>
<wire>
<ID>2583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-781,-4731,-781,-4723.5</points>
<connection>
<GID>2411</GID>
<name>IN_0</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-784.5,-4723.5,-781,-4723.5</points>
<connection>
<GID>2405</GID>
<name>OUT_0</name></connection>
<intersection>-781 0</intersection></hsegment></shape></wire>
<wire>
<ID>2584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-768,-4730.5,-768,-4723.5</points>
<connection>
<GID>2412</GID>
<name>IN_0</name></connection>
<intersection>-4723.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-771.5,-4723.5,-768,-4723.5</points>
<connection>
<GID>2406</GID>
<name>OUT_0</name></connection>
<intersection>-768 0</intersection></hsegment></shape></wire>
<wire>
<ID>2585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-835.5,-4740.5,-835.5,-4735</points>
<connection>
<GID>2407</GID>
<name>OUT_0</name></connection>
<intersection>-4740.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-820.5,-4746.5,-820.5,-4740.5</points>
<connection>
<GID>2413</GID>
<name>IN_3</name></connection>
<intersection>-4740.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-835.5,-4740.5,-820.5,-4740.5</points>
<intersection>-835.5 0</intersection>
<intersection>-820.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-820.5,-4740,-820.5,-4735</points>
<connection>
<GID>2408</GID>
<name>OUT_0</name></connection>
<intersection>-4740 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-818.5,-4746.5,-818.5,-4740</points>
<connection>
<GID>2413</GID>
<name>IN_2</name></connection>
<intersection>-4740 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-820.5,-4740,-818.5,-4740</points>
<intersection>-820.5 0</intersection>
<intersection>-818.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805.5,-4740.5,-805.5,-4735</points>
<connection>
<GID>2409</GID>
<name>OUT_0</name></connection>
<intersection>-4740.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-816.5,-4746.5,-816.5,-4740.5</points>
<connection>
<GID>2413</GID>
<name>IN_1</name></connection>
<intersection>-4740.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-816.5,-4740.5,-805.5,-4740.5</points>
<intersection>-816.5 1</intersection>
<intersection>-805.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-794,-4741.5,-794,-4734.5</points>
<connection>
<GID>2410</GID>
<name>OUT_0</name></connection>
<intersection>-4741.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-814.5,-4746.5,-814.5,-4741.5</points>
<connection>
<GID>2413</GID>
<name>IN_0</name></connection>
<intersection>-4741.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-814.5,-4741.5,-794,-4741.5</points>
<intersection>-814.5 1</intersection>
<intersection>-794 0</intersection></hsegment></shape></wire>
<wire>
<ID>2589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-781,-4740,-781,-4735</points>
<connection>
<GID>2411</GID>
<name>OUT_0</name></connection>
<intersection>-4740 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-782,-4745.5,-782,-4740</points>
<connection>
<GID>2415</GID>
<name>IN_1</name></connection>
<intersection>-4740 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-782,-4740,-781,-4740</points>
<intersection>-782 1</intersection>
<intersection>-781 0</intersection></hsegment></shape></wire>
<wire>
<ID>2590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-768,-4740,-768,-4734.5</points>
<connection>
<GID>2412</GID>
<name>OUT_0</name></connection>
<intersection>-4740 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-780,-4745.5,-780,-4740</points>
<connection>
<GID>2415</GID>
<name>IN_0</name></connection>
<intersection>-4740 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-780,-4740,-768,-4740</points>
<intersection>-780 1</intersection>
<intersection>-768 0</intersection></hsegment></shape></wire>
<wire>
<ID>2591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-817.5,-4755.5,-817.5,-4752.5</points>
<connection>
<GID>2413</GID>
<name>OUT</name></connection>
<intersection>-4755.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-804.5,-4768.5,-804.5,-4755.5</points>
<connection>
<GID>2416</GID>
<name>IN_1</name></connection>
<intersection>-4763.5 7</intersection>
<intersection>-4755.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-868,-4755.5,-804.5,-4755.5</points>
<connection>
<GID>1977</GID>
<name>IN_0</name></connection>
<intersection>-817.5 0</intersection>
<intersection>-804.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-804.5,-4763.5,-793,-4763.5</points>
<connection>
<GID>2429</GID>
<name>IN_0</name></connection>
<intersection>-804.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-781,-4755,-781,-4751.5</points>
<connection>
<GID>2415</GID>
<name>OUT</name></connection>
<intersection>-4755 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-802.5,-4768.5,-802.5,-4755</points>
<connection>
<GID>2416</GID>
<name>IN_0</name></connection>
<intersection>-4765.5 6</intersection>
<intersection>-4757.5 7</intersection>
<intersection>-4755 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-802.5,-4755,-781,-4755</points>
<intersection>-802.5 1</intersection>
<intersection>-781 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-802.5,-4765.5,-793,-4765.5</points>
<connection>
<GID>2429</GID>
<name>IN_1</name></connection>
<intersection>-802.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-908.5,-4757.5,-802.5,-4757.5</points>
<connection>
<GID>1967</GID>
<name>IN_0</name></connection>
<intersection>-802.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-929.5,-4677.5,-870.5,-4677.5</points>
<connection>
<GID>2434</GID>
<name>OUT</name></connection>
<connection>
<GID>2426</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-847.5,-4713.5,-847.5,-4677.5</points>
<connection>
<GID>2417</GID>
<name>IN_1</name></connection>
<intersection>-4677.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-864.5,-4677.5,-847.5,-4677.5</points>
<connection>
<GID>2426</GID>
<name>Q</name></connection>
<intersection>-847.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-930,-4667.5,-883.5,-4667.5</points>
<connection>
<GID>2435</GID>
<name>OUT</name></connection>
<connection>
<GID>2427</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-834,-4713.5,-834,-4667.5</points>
<connection>
<GID>2418</GID>
<name>IN_1</name></connection>
<intersection>-4667.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-877.5,-4667.5,-834,-4667.5</points>
<connection>
<GID>2427</GID>
<name>Q</name></connection>
<intersection>-834 0</intersection></hsegment></shape></wire>
<wire>
<ID>2597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-931.5,-4656.5,-896.5,-4656.5</points>
<connection>
<GID>2436</GID>
<name>OUT</name></connection>
<connection>
<GID>2428</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-821,-4713.5,-821,-4656.5</points>
<connection>
<GID>2419</GID>
<name>IN_1</name></connection>
<intersection>-4656.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-890.5,-4656.5,-821,-4656.5</points>
<connection>
<GID>2428</GID>
<name>Q</name></connection>
<intersection>-821 0</intersection></hsegment></shape></wire>
<wire>
<ID>2599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-932,-4647.5,-904,-4647.5</points>
<connection>
<GID>2437</GID>
<name>OUT</name></connection>
<connection>
<GID>2430</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808,-4713.5,-808,-4647.5</points>
<connection>
<GID>2420</GID>
<name>IN_1</name></connection>
<intersection>-4647.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-898,-4647.5,-808,-4647.5</points>
<connection>
<GID>2430</GID>
<name>Q</name></connection>
<intersection>-808 0</intersection></hsegment></shape></wire>
<wire>
<ID>2601</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-933,-4640,-912.5,-4640</points>
<connection>
<GID>2438</GID>
<name>OUT</name></connection>
<connection>
<GID>2431</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795.5,-4714,-795.5,-4640</points>
<connection>
<GID>2421</GID>
<name>IN_1</name></connection>
<intersection>-4640 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-906.5,-4640,-795.5,-4640</points>
<connection>
<GID>2431</GID>
<name>Q</name></connection>
<intersection>-795.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2603</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-934,-4632.5,-921.5,-4632.5</points>
<connection>
<GID>2439</GID>
<name>OUT</name></connection>
<connection>
<GID>2432</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-783,-4714,-783,-4632.5</points>
<connection>
<GID>2423</GID>
<name>IN_1</name></connection>
<intersection>-4632.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-915.5,-4632.5,-783,-4632.5</points>
<connection>
<GID>2432</GID>
<name>Q</name></connection>
<intersection>-783 0</intersection></hsegment></shape></wire>
<wire>
<ID>2605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-926.5,-4679.5,-926.5,-4628.5</points>
<connection>
<GID>2433</GID>
<name>OUT_0</name></connection>
<intersection>-4679.5 7</intersection>
<intersection>-4669.5 5</intersection>
<intersection>-4658.5 8</intersection>
<intersection>-4649.5 3</intersection>
<intersection>-4642 9</intersection>
<intersection>-4634.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-926.5,-4634.5,-921.5,-4634.5</points>
<connection>
<GID>2432</GID>
<name>clock</name></connection>
<intersection>-926.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-926.5,-4649.5,-904,-4649.5</points>
<connection>
<GID>2430</GID>
<name>clock</name></connection>
<intersection>-926.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-926.5,-4669.5,-883.5,-4669.5</points>
<connection>
<GID>2427</GID>
<name>clock</name></connection>
<intersection>-926.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-926.5,-4679.5,-870.5,-4679.5</points>
<connection>
<GID>2426</GID>
<name>clock</name></connection>
<intersection>-926.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-926.5,-4658.5,-896.5,-4658.5</points>
<connection>
<GID>2428</GID>
<name>clock</name></connection>
<intersection>-926.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-926.5,-4642,-912.5,-4642</points>
<connection>
<GID>2431</GID>
<name>clock</name></connection>
<intersection>-926.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-957.5,-4993.5,-957.5,-4825</points>
<intersection>-4993.5 13</intersection>
<intersection>-4903.5 1</intersection>
<intersection>-4893.5 3</intersection>
<intersection>-4882.5 5</intersection>
<intersection>-4873.5 7</intersection>
<intersection>-4866 9</intersection>
<intersection>-4832.5 11</intersection>
<intersection>-4825 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-957.5,-4903.5,-926.5,-4903.5</points>
<connection>
<GID>2472</GID>
<name>IN_0</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-957.5,-4893.5,-927,-4893.5</points>
<connection>
<GID>2473</GID>
<name>IN_0</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-957.5,-4882.5,-928.5,-4882.5</points>
<connection>
<GID>2474</GID>
<name>IN_0</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-957.5,-4873.5,-929,-4873.5</points>
<connection>
<GID>2475</GID>
<name>IN_0</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-957.5,-4866,-930,-4866</points>
<connection>
<GID>2476</GID>
<name>IN_0</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-957.5,-4832.5,-775,-4832.5</points>
<intersection>-957.5 0</intersection>
<intersection>-931 15</intersection>
<intersection>-775 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-957.5,-4993.5,-772,-4993.5</points>
<connection>
<GID>1893</GID>
<name>IN_1</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-775,-4832.5,-775,-4790</points>
<connection>
<GID>2057</GID>
<name>IN_1</name></connection>
<intersection>-4832.5 11</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-931,-4858.5,-931,-4832.5</points>
<connection>
<GID>2477</GID>
<name>IN_0</name></connection>
<intersection>-4832.5 11</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-959.5,-4825,-957.5,-4825</points>
<connection>
<GID>2130</GID>
<name>OUT</name></connection>
<intersection>-957.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-837.5,-4950,-837.5,-4946.5</points>
<connection>
<GID>2456</GID>
<name>OUT</name></connection>
<intersection>-4950 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-837.5,-4950,-836.5,-4950</points>
<connection>
<GID>2478</GID>
<name>IN_0</name></connection>
<intersection>-837.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-824,-4950.5,-824,-4946.5</points>
<connection>
<GID>2457</GID>
<name>OUT</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-824,-4950.5,-820.5,-4950.5</points>
<connection>
<GID>2441</GID>
<name>IN_0</name></connection>
<intersection>-824 0</intersection></hsegment></shape></wire>
<wire>
<ID>2609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-811,-4950.5,-811,-4946.5</points>
<connection>
<GID>2458</GID>
<name>OUT</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-811,-4950.5,-807,-4950.5</points>
<connection>
<GID>2442</GID>
<name>IN_0</name></connection>
<intersection>-811 0</intersection></hsegment></shape></wire>
<wire>
<ID>2610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795,-4950.5,-795,-4946.5</points>
<intersection>-4950.5 1</intersection>
<intersection>-4946.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-795,-4950.5,-792,-4950.5</points>
<connection>
<GID>2443</GID>
<name>IN_0</name></connection>
<intersection>-795 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-798,-4946.5,-795,-4946.5</points>
<connection>
<GID>2459</GID>
<name>OUT</name></connection>
<intersection>-795 0</intersection></hsegment></shape></wire>
<wire>
<ID>2611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-785.5,-4949,-785.5,-4947</points>
<connection>
<GID>2460</GID>
<name>OUT</name></connection>
<intersection>-4949 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-785.5,-4949,-781.5,-4949</points>
<intersection>-785.5 0</intersection>
<intersection>-781.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-781.5,-4950.5,-781.5,-4949</points>
<connection>
<GID>2444</GID>
<name>IN_0</name></connection>
<intersection>-4949 1</intersection></vsegment></shape></wire>
<wire>
<ID>2612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-773,-4949,-773,-4947</points>
<connection>
<GID>2461</GID>
<name>OUT</name></connection>
<intersection>-4949 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-773,-4949,-768.5,-4949</points>
<intersection>-773 0</intersection>
<intersection>-768.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-768.5,-4950.5,-768.5,-4949</points>
<connection>
<GID>2445</GID>
<name>IN_0</name></connection>
<intersection>-4949 1</intersection></vsegment></shape></wire>
<wire>
<ID>2613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-826.5,-4958,-826.5,-4950</points>
<connection>
<GID>2446</GID>
<name>IN_0</name></connection>
<intersection>-4950 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-830.5,-4950,-826.5,-4950</points>
<connection>
<GID>2478</GID>
<name>OUT_0</name></connection>
<intersection>-826.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-811.5,-4958,-811.5,-4950.5</points>
<connection>
<GID>2447</GID>
<name>IN_0</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-814.5,-4950.5,-811.5,-4950.5</points>
<connection>
<GID>2441</GID>
<name>OUT_0</name></connection>
<intersection>-811.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-796.5,-4958,-796.5,-4950.5</points>
<connection>
<GID>2448</GID>
<name>IN_0</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-801,-4950.5,-796.5,-4950.5</points>
<connection>
<GID>2442</GID>
<name>OUT_0</name></connection>
<intersection>-796.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-785,-4957.5,-785,-4950.5</points>
<connection>
<GID>2449</GID>
<name>IN_0</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-786,-4950.5,-785,-4950.5</points>
<connection>
<GID>2443</GID>
<name>OUT_0</name></connection>
<intersection>-785 0</intersection></hsegment></shape></wire>
<wire>
<ID>2617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-772,-4958,-772,-4950.5</points>
<connection>
<GID>2450</GID>
<name>IN_0</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-775.5,-4950.5,-772,-4950.5</points>
<connection>
<GID>2444</GID>
<name>OUT_0</name></connection>
<intersection>-772 0</intersection></hsegment></shape></wire>
<wire>
<ID>2618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-759,-4957.5,-759,-4950.5</points>
<connection>
<GID>2451</GID>
<name>IN_0</name></connection>
<intersection>-4950.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-762.5,-4950.5,-759,-4950.5</points>
<connection>
<GID>2445</GID>
<name>OUT_0</name></connection>
<intersection>-759 0</intersection></hsegment></shape></wire>
<wire>
<ID>2619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-826.5,-4967.5,-826.5,-4962</points>
<connection>
<GID>2446</GID>
<name>OUT_0</name></connection>
<intersection>-4967.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-811.5,-4973.5,-811.5,-4967.5</points>
<connection>
<GID>2452</GID>
<name>IN_3</name></connection>
<intersection>-4967.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-826.5,-4967.5,-811.5,-4967.5</points>
<intersection>-826.5 0</intersection>
<intersection>-811.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-811.5,-4967,-811.5,-4962</points>
<connection>
<GID>2447</GID>
<name>OUT_0</name></connection>
<intersection>-4967 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-809.5,-4973.5,-809.5,-4967</points>
<connection>
<GID>2452</GID>
<name>IN_2</name></connection>
<intersection>-4967 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-811.5,-4967,-809.5,-4967</points>
<intersection>-811.5 0</intersection>
<intersection>-809.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-796.5,-4967.5,-796.5,-4962</points>
<connection>
<GID>2448</GID>
<name>OUT_0</name></connection>
<intersection>-4967.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-807.5,-4973.5,-807.5,-4967.5</points>
<connection>
<GID>2452</GID>
<name>IN_1</name></connection>
<intersection>-4967.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-807.5,-4967.5,-796.5,-4967.5</points>
<intersection>-807.5 1</intersection>
<intersection>-796.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-785,-4968.5,-785,-4961.5</points>
<connection>
<GID>2449</GID>
<name>OUT_0</name></connection>
<intersection>-4968.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-805.5,-4973.5,-805.5,-4968.5</points>
<connection>
<GID>2452</GID>
<name>IN_0</name></connection>
<intersection>-4968.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-805.5,-4968.5,-785,-4968.5</points>
<intersection>-805.5 1</intersection>
<intersection>-785 0</intersection></hsegment></shape></wire>
<wire>
<ID>2623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-772,-4967,-772,-4962</points>
<connection>
<GID>2450</GID>
<name>OUT_0</name></connection>
<intersection>-4967 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-773,-4972.5,-773,-4967</points>
<connection>
<GID>2454</GID>
<name>IN_1</name></connection>
<intersection>-4967 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-773,-4967,-772,-4967</points>
<intersection>-773 1</intersection>
<intersection>-772 0</intersection></hsegment></shape></wire>
<wire>
<ID>2624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-759,-4967,-759,-4961.5</points>
<connection>
<GID>2451</GID>
<name>OUT_0</name></connection>
<intersection>-4967 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-771,-4972.5,-771,-4967</points>
<connection>
<GID>2454</GID>
<name>IN_0</name></connection>
<intersection>-4967 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-771,-4967,-759,-4967</points>
<intersection>-771 1</intersection>
<intersection>-759 0</intersection></hsegment></shape></wire>
<wire>
<ID>2625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808.5,-4984,-808.5,-4979.5</points>
<connection>
<GID>2452</GID>
<name>OUT</name></connection>
<intersection>-4984 8</intersection>
<intersection>-4982.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-795.5,-4995.5,-795.5,-4982.5</points>
<connection>
<GID>2455</GID>
<name>IN_1</name></connection>
<intersection>-4990.5 7</intersection>
<intersection>-4982.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-808.5,-4982.5,-795.5,-4982.5</points>
<intersection>-808.5 0</intersection>
<intersection>-795.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-795.5,-4990.5,-784,-4990.5</points>
<connection>
<GID>2467</GID>
<name>IN_0</name></connection>
<intersection>-795.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-845.5,-4984,-808.5,-4984</points>
<connection>
<GID>1988</GID>
<name>IN_0</name></connection>
<intersection>-808.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-772,-4982,-772,-4978.5</points>
<connection>
<GID>2454</GID>
<name>OUT</name></connection>
<intersection>-4982 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-793.5,-4995.5,-793.5,-4982</points>
<connection>
<GID>2455</GID>
<name>IN_0</name></connection>
<intersection>-4992.5 6</intersection>
<intersection>-4986 7</intersection>
<intersection>-4982 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-793.5,-4982,-772,-4982</points>
<intersection>-793.5 1</intersection>
<intersection>-772 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-793.5,-4992.5,-784,-4992.5</points>
<connection>
<GID>2467</GID>
<name>IN_1</name></connection>
<intersection>-793.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-886,-4986,-793.5,-4986</points>
<connection>
<GID>1981</GID>
<name>IN_0</name></connection>
<intersection>-793.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-920.5,-4904.5,-861.5,-4904.5</points>
<connection>
<GID>2472</GID>
<name>OUT</name></connection>
<connection>
<GID>2464</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-838.5,-4940.5,-838.5,-4904.5</points>
<connection>
<GID>2456</GID>
<name>IN_1</name></connection>
<intersection>-4904.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-855.5,-4904.5,-838.5,-4904.5</points>
<connection>
<GID>2464</GID>
<name>Q</name></connection>
<intersection>-838.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-921,-4894.5,-874.5,-4894.5</points>
<connection>
<GID>2473</GID>
<name>OUT</name></connection>
<connection>
<GID>2465</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-825,-4940.5,-825,-4894.5</points>
<connection>
<GID>2457</GID>
<name>IN_1</name></connection>
<intersection>-4894.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-868.5,-4894.5,-825,-4894.5</points>
<connection>
<GID>2465</GID>
<name>Q</name></connection>
<intersection>-825 0</intersection></hsegment></shape></wire>
<wire>
<ID>2631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-922.5,-4883.5,-887.5,-4883.5</points>
<connection>
<GID>2474</GID>
<name>OUT</name></connection>
<connection>
<GID>2466</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-812,-4940.5,-812,-4883.5</points>
<connection>
<GID>2458</GID>
<name>IN_1</name></connection>
<intersection>-4883.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-881.5,-4883.5,-812,-4883.5</points>
<connection>
<GID>2466</GID>
<name>Q</name></connection>
<intersection>-812 0</intersection></hsegment></shape></wire>
<wire>
<ID>2633</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-923,-4874.5,-895,-4874.5</points>
<connection>
<GID>2475</GID>
<name>OUT</name></connection>
<connection>
<GID>2468</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-799,-4940.5,-799,-4874.5</points>
<connection>
<GID>2459</GID>
<name>IN_1</name></connection>
<intersection>-4874.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-889,-4874.5,-799,-4874.5</points>
<connection>
<GID>2468</GID>
<name>Q</name></connection>
<intersection>-799 0</intersection></hsegment></shape></wire>
<wire>
<ID>2635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-924,-4867,-903.5,-4867</points>
<connection>
<GID>2476</GID>
<name>OUT</name></connection>
<connection>
<GID>2469</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-786.5,-4941,-786.5,-4867</points>
<connection>
<GID>2460</GID>
<name>IN_1</name></connection>
<intersection>-4867 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-897.5,-4867,-786.5,-4867</points>
<connection>
<GID>2469</GID>
<name>Q</name></connection>
<intersection>-786.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-925,-4859.5,-912.5,-4859.5</points>
<connection>
<GID>2477</GID>
<name>OUT</name></connection>
<connection>
<GID>2470</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-774,-4941,-774,-4859.5</points>
<connection>
<GID>2461</GID>
<name>IN_1</name></connection>
<intersection>-4859.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-906.5,-4859.5,-774,-4859.5</points>
<connection>
<GID>2470</GID>
<name>Q</name></connection>
<intersection>-774 0</intersection></hsegment></shape></wire>
<wire>
<ID>2639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-917.5,-4906.5,-917.5,-4855.5</points>
<connection>
<GID>2471</GID>
<name>OUT_0</name></connection>
<intersection>-4906.5 7</intersection>
<intersection>-4896.5 5</intersection>
<intersection>-4885.5 8</intersection>
<intersection>-4876.5 3</intersection>
<intersection>-4869 9</intersection>
<intersection>-4861.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-917.5,-4861.5,-912.5,-4861.5</points>
<connection>
<GID>2470</GID>
<name>clock</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-917.5,-4876.5,-895,-4876.5</points>
<connection>
<GID>2468</GID>
<name>clock</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-917.5,-4896.5,-874.5,-4896.5</points>
<connection>
<GID>2465</GID>
<name>clock</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-917.5,-4906.5,-861.5,-4906.5</points>
<connection>
<GID>2464</GID>
<name>clock</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-917.5,-4885.5,-887.5,-4885.5</points>
<connection>
<GID>2466</GID>
<name>clock</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-917.5,-4869,-903.5,-4869</points>
<connection>
<GID>2469</GID>
<name>clock</name></connection>
<intersection>-917.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-871.5,-3714.5,-871.5,-3710</points>
<connection>
<GID>2162</GID>
<name>IN_1</name></connection>
<intersection>-3710 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-898,-3710,-871.5,-3710</points>
<connection>
<GID>2368</GID>
<name>Q</name></connection>
<intersection>-871.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2641</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-956.5,-3701.5,-912,-3701.5</points>
<connection>
<GID>2347</GID>
<name>OUT</name></connection>
<connection>
<GID>2370</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-858,-3714.5,-858,-3701.5</points>
<connection>
<GID>2163</GID>
<name>IN_1</name></connection>
<intersection>-3701.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-906,-3701.5,-858,-3701.5</points>
<connection>
<GID>2370</GID>
<name>Q</name></connection>
<intersection>-858 0</intersection></hsegment></shape></wire>
<wire>
<ID>2643</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-957,-3693,-919,-3693</points>
<connection>
<GID>2348</GID>
<name>OUT</name></connection>
<connection>
<GID>2371</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-845,-3714.5,-845,-3693</points>
<connection>
<GID>2164</GID>
<name>IN_1</name></connection>
<intersection>-3693 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-913,-3693,-845,-3693</points>
<connection>
<GID>2371</GID>
<name>Q</name></connection>
<intersection>-845 0</intersection></hsegment></shape></wire>
<wire>
<ID>2645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-957.5,-3685,-928,-3685</points>
<connection>
<GID>2349</GID>
<name>OUT</name></connection>
<connection>
<GID>2372</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-832,-3714.5,-832,-3685</points>
<connection>
<GID>2165</GID>
<name>IN_1</name></connection>
<intersection>-3685 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-922,-3685,-832,-3685</points>
<connection>
<GID>2372</GID>
<name>Q</name></connection>
<intersection>-832 0</intersection></hsegment></shape></wire>
<wire>
<ID>2647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-958,-3676.5,-935,-3676.5</points>
<connection>
<GID>2350</GID>
<name>OUT</name></connection>
<connection>
<GID>2374</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-819.5,-3715,-819.5,-3676.5</points>
<connection>
<GID>2166</GID>
<name>IN_1</name></connection>
<intersection>-3676.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-929,-3676.5,-819.5,-3676.5</points>
<connection>
<GID>2374</GID>
<name>Q</name></connection>
<intersection>-819.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2649</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-958,-3668,-943,-3668</points>
<connection>
<GID>2351</GID>
<name>OUT</name></connection>
<connection>
<GID>2375</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-807,-3715,-807,-3668</points>
<connection>
<GID>2167</GID>
<name>IN_1</name></connection>
<intersection>-3668 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-937,-3668,-807,-3668</points>
<connection>
<GID>2375</GID>
<name>Q</name></connection>
<intersection>-807 0</intersection></hsegment></shape></wire>
<wire>
<ID>2651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-948,-3712,-948,-3660</points>
<connection>
<GID>2387</GID>
<name>OUT_0</name></connection>
<intersection>-3712 7</intersection>
<intersection>-3703.5 5</intersection>
<intersection>-3695 8</intersection>
<intersection>-3687 3</intersection>
<intersection>-3678.5 9</intersection>
<intersection>-3670 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-948,-3670,-943,-3670</points>
<connection>
<GID>2375</GID>
<name>clock</name></connection>
<intersection>-948 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-948,-3687,-928,-3687</points>
<connection>
<GID>2372</GID>
<name>clock</name></connection>
<intersection>-948 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-948,-3703.5,-912,-3703.5</points>
<connection>
<GID>2370</GID>
<name>clock</name></connection>
<intersection>-948 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-948,-3712,-904,-3712</points>
<connection>
<GID>2368</GID>
<name>clock</name></connection>
<intersection>-948 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-948,-3695,-919,-3695</points>
<connection>
<GID>2371</GID>
<name>clock</name></connection>
<intersection>-948 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-948,-3678.5,-935,-3678.5</points>
<connection>
<GID>2374</GID>
<name>clock</name></connection>
<intersection>-948 0</intersection></hsegment></shape></wire>
<wire>
<ID>2652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-950.5,-3555.5,-950.5,-3504.5</points>
<connection>
<GID>2391</GID>
<name>OUT_0</name></connection>
<intersection>-3555.5 7</intersection>
<intersection>-3545.5 5</intersection>
<intersection>-3534.5 8</intersection>
<intersection>-3525.5 3</intersection>
<intersection>-3518 9</intersection>
<intersection>-3510.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-950.5,-3510.5,-945,-3510.5</points>
<connection>
<GID>2367</GID>
<name>clock</name></connection>
<intersection>-950.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-950.5,-3525.5,-927.5,-3525.5</points>
<connection>
<GID>2365</GID>
<name>clock</name></connection>
<intersection>-950.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-950.5,-3545.5,-907,-3545.5</points>
<connection>
<GID>2363</GID>
<name>clock</name></connection>
<intersection>-950.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-950.5,-3555.5,-894,-3555.5</points>
<connection>
<GID>2360</GID>
<name>clock</name></connection>
<intersection>-950.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-950.5,-3534.5,-920,-3534.5</points>
<connection>
<GID>2364</GID>
<name>clock</name></connection>
<intersection>-950.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-950.5,-3518,-936,-3518</points>
<connection>
<GID>2366</GID>
<name>clock</name></connection>
<intersection>-950.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-725,-3721.5,-725,-3487</points>
<intersection>-3721.5 17</intersection>
<intersection>-3559.5 3</intersection>
<intersection>-3487 26</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-942,-3559.5,-725,-3559.5</points>
<connection>
<GID>2360</GID>
<name>clear</name></connection>
<intersection>-942 27</intersection>
<intersection>-933 28</intersection>
<intersection>-924.5 29</intersection>
<intersection>-917 30</intersection>
<intersection>-904 31</intersection>
<intersection>-725 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-940,-3721.5,-725,-3721.5</points>
<intersection>-940 33</intersection>
<intersection>-932 34</intersection>
<intersection>-925 35</intersection>
<intersection>-916 36</intersection>
<intersection>-909 37</intersection>
<intersection>-901 38</intersection>
<intersection>-725.5 39</intersection>
<intersection>-725 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-787.5,-3487,-725,-3487</points>
<intersection>-787.5 32</intersection>
<intersection>-725 0</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>-942,-3559.5,-942,-3514.5</points>
<connection>
<GID>2367</GID>
<name>clear</name></connection>
<intersection>-3559.5 3</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-933,-3559.5,-933,-3522</points>
<connection>
<GID>2366</GID>
<name>clear</name></connection>
<intersection>-3559.5 3</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>-924.5,-3559.5,-924.5,-3529.5</points>
<connection>
<GID>2365</GID>
<name>clear</name></connection>
<intersection>-3559.5 3</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-917,-3559.5,-917,-3538.5</points>
<connection>
<GID>2364</GID>
<name>clear</name></connection>
<intersection>-3559.5 3</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-904,-3559.5,-904,-3549.5</points>
<connection>
<GID>2363</GID>
<name>clear</name></connection>
<intersection>-3559.5 3</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-787.5,-3487,-787.5,-3480.5</points>
<connection>
<GID>2395</GID>
<name>OUT_0</name></connection>
<intersection>-3487 26</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>-940,-3721.5,-940,-3674</points>
<connection>
<GID>2375</GID>
<name>clear</name></connection>
<intersection>-3721.5 17</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-932,-3721.5,-932,-3682.5</points>
<connection>
<GID>2374</GID>
<name>clear</name></connection>
<intersection>-3721.5 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>-925,-3721.5,-925,-3691</points>
<connection>
<GID>2372</GID>
<name>clear</name></connection>
<intersection>-3721.5 17</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>-916,-3721.5,-916,-3699</points>
<connection>
<GID>2371</GID>
<name>clear</name></connection>
<intersection>-3721.5 17</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>-909,-3721.5,-909,-3707.5</points>
<connection>
<GID>2370</GID>
<name>clear</name></connection>
<intersection>-3721.5 17</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>-901,-3721.5,-901,-3716</points>
<connection>
<GID>2368</GID>
<name>clear</name></connection>
<intersection>-3721.5 17</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>-725.5,-4449.5,-725.5,-3721.5</points>
<intersection>-4449.5 105</intersection>
<intersection>-4227.5 84</intersection>
<intersection>-4036 64</intersection>
<intersection>-3852.5 43</intersection>
<intersection>-3721.5 17</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>-933,-3852.5,-725.5,-3852.5</points>
<intersection>-933 53</intersection>
<intersection>-923.5 54</intersection>
<intersection>-915 55</intersection>
<intersection>-907.5 56</intersection>
<intersection>-894.5 57</intersection>
<intersection>-881.5 59</intersection>
<intersection>-725.5 39</intersection></hsegment>
<vsegment>
<ID>53</ID>
<points>-933,-3852.5,-933,-3801.5</points>
<intersection>-3852.5 43</intersection>
<intersection>-3801.5 58</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>-923.5,-3852.5,-923.5,-3809</points>
<connection>
<GID>1945</GID>
<name>clear</name></connection>
<intersection>-3852.5 43</intersection></vsegment>
<vsegment>
<ID>55</ID>
<points>-915,-3852.5,-915,-3816.5</points>
<connection>
<GID>1944</GID>
<name>clear</name></connection>
<intersection>-3852.5 43</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>-907.5,-3852.5,-907.5,-3825.5</points>
<connection>
<GID>1942</GID>
<name>clear</name></connection>
<intersection>-3852.5 43</intersection></vsegment>
<vsegment>
<ID>57</ID>
<points>-894.5,-3852.5,-894.5,-3836.5</points>
<connection>
<GID>1941</GID>
<name>clear</name></connection>
<intersection>-3852.5 43</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>-933,-3801.5,-932.5,-3801.5</points>
<connection>
<GID>1947</GID>
<name>clear</name></connection>
<intersection>-933 53</intersection></hsegment>
<vsegment>
<ID>59</ID>
<points>-881.5,-3852.5,-881.5,-3846.5</points>
<connection>
<GID>1940</GID>
<name>clear</name></connection>
<intersection>-3852.5 43</intersection></vsegment>
<hsegment>
<ID>64</ID>
<points>-924.5,-4036,-725.5,-4036</points>
<intersection>-924.5 74</intersection>
<intersection>-915.5 75</intersection>
<intersection>-907 76</intersection>
<intersection>-899.5 77</intersection>
<intersection>-886.5 78</intersection>
<intersection>-873.5 79</intersection>
<intersection>-725.5 39</intersection></hsegment>
<vsegment>
<ID>74</ID>
<points>-924.5,-4036,-924.5,-3983.5</points>
<connection>
<GID>2023</GID>
<name>clear</name></connection>
<intersection>-4036 64</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>-915.5,-4036,-915.5,-3991</points>
<connection>
<GID>2022</GID>
<name>clear</name></connection>
<intersection>-4036 64</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>-907,-4036,-907,-3998.5</points>
<connection>
<GID>2021</GID>
<name>clear</name></connection>
<intersection>-4036 64</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>-899.5,-4036,-899.5,-4007.5</points>
<connection>
<GID>2019</GID>
<name>clear</name></connection>
<intersection>-4036 64</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>-886.5,-4036,-886.5,-4018.5</points>
<connection>
<GID>2018</GID>
<name>clear</name></connection>
<intersection>-4036 64</intersection></vsegment>
<vsegment>
<ID>79</ID>
<points>-873.5,-4036,-873.5,-4028.5</points>
<connection>
<GID>2017</GID>
<name>clear</name></connection>
<intersection>-4036 64</intersection></vsegment>
<hsegment>
<ID>84</ID>
<points>-914,-4227.5,-725.5,-4227.5</points>
<connection>
<GID>2127</GID>
<name>clear</name></connection>
<intersection>-914 94</intersection>
<intersection>-905 95</intersection>
<intersection>-896.5 100</intersection>
<intersection>-889 97</intersection>
<intersection>-876 98</intersection>
<intersection>-725.5 39</intersection></hsegment>
<vsegment>
<ID>94</ID>
<points>-914,-4227.5,-914,-4182.5</points>
<connection>
<GID>2138</GID>
<name>clear</name></connection>
<intersection>-4227.5 84</intersection></vsegment>
<vsegment>
<ID>95</ID>
<points>-905,-4227.5,-905,-4190</points>
<connection>
<GID>2137</GID>
<name>clear</name></connection>
<intersection>-4227.5 84</intersection></vsegment>
<vsegment>
<ID>97</ID>
<points>-889,-4227.5,-889,-4206.5</points>
<connection>
<GID>2131</GID>
<name>clear</name></connection>
<intersection>-4227.5 84</intersection></vsegment>
<vsegment>
<ID>98</ID>
<points>-876,-4227.5,-876,-4217.5</points>
<connection>
<GID>2129</GID>
<name>clear</name></connection>
<intersection>-4227.5 84</intersection></vsegment>
<vsegment>
<ID>100</ID>
<points>-896.5,-4227.5,-896.5,-4197.5</points>
<connection>
<GID>2135</GID>
<name>clear</name></connection>
<intersection>-4227.5 84</intersection></vsegment>
<hsegment>
<ID>105</ID>
<points>-920.5,-4449.5,-725.5,-4449.5</points>
<connection>
<GID>2377</GID>
<name>clear</name></connection>
<intersection>-920.5 115</intersection>
<intersection>-911.5 116</intersection>
<intersection>-903 117</intersection>
<intersection>-895.5 118</intersection>
<intersection>-882.5 119</intersection>
<intersection>-726 120</intersection>
<intersection>-725.5 39</intersection></hsegment>
<vsegment>
<ID>115</ID>
<points>-920.5,-4449.5,-920.5,-4404.5</points>
<connection>
<GID>2389</GID>
<name>clear</name></connection>
<intersection>-4449.5 105</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>-911.5,-4449.5,-911.5,-4412</points>
<connection>
<GID>2386</GID>
<name>clear</name></connection>
<intersection>-4449.5 105</intersection></vsegment>
<vsegment>
<ID>117</ID>
<points>-903,-4449.5,-903,-4419.5</points>
<connection>
<GID>2384</GID>
<name>clear</name></connection>
<intersection>-4449.5 105</intersection></vsegment>
<vsegment>
<ID>118</ID>
<points>-895.5,-4449.5,-895.5,-4428.5</points>
<connection>
<GID>2380</GID>
<name>clear</name></connection>
<intersection>-4449.5 105</intersection></vsegment>
<vsegment>
<ID>119</ID>
<points>-882.5,-4449.5,-882.5,-4439.5</points>
<connection>
<GID>2379</GID>
<name>clear</name></connection>
<intersection>-4449.5 105</intersection></vsegment>
<vsegment>
<ID>120</ID>
<points>-726,-4683.5,-726,-4449.5</points>
<intersection>-4683.5 124</intersection>
<intersection>-4449.5 105</intersection></vsegment>
<hsegment>
<ID>124</ID>
<points>-918.5,-4683.5,-726,-4683.5</points>
<connection>
<GID>2426</GID>
<name>clear</name></connection>
<intersection>-918.5 134</intersection>
<intersection>-909.5 135</intersection>
<intersection>-901 136</intersection>
<intersection>-893.5 137</intersection>
<intersection>-880.5 138</intersection>
<intersection>-726.5 139</intersection>
<intersection>-726 120</intersection></hsegment>
<vsegment>
<ID>134</ID>
<points>-918.5,-4683.5,-918.5,-4638.5</points>
<connection>
<GID>2432</GID>
<name>clear</name></connection>
<intersection>-4683.5 124</intersection></vsegment>
<vsegment>
<ID>135</ID>
<points>-909.5,-4683.5,-909.5,-4646</points>
<connection>
<GID>2431</GID>
<name>clear</name></connection>
<intersection>-4683.5 124</intersection></vsegment>
<vsegment>
<ID>136</ID>
<points>-901,-4683.5,-901,-4653.5</points>
<connection>
<GID>2430</GID>
<name>clear</name></connection>
<intersection>-4683.5 124</intersection></vsegment>
<vsegment>
<ID>137</ID>
<points>-893.5,-4683.5,-893.5,-4662.5</points>
<connection>
<GID>2428</GID>
<name>clear</name></connection>
<intersection>-4683.5 124</intersection></vsegment>
<vsegment>
<ID>138</ID>
<points>-880.5,-4683.5,-880.5,-4673.5</points>
<connection>
<GID>2427</GID>
<name>clear</name></connection>
<intersection>-4683.5 124</intersection></vsegment>
<vsegment>
<ID>139</ID>
<points>-726.5,-4910.5,-726.5,-4683.5</points>
<intersection>-4910.5 143</intersection>
<intersection>-4683.5 124</intersection></vsegment>
<hsegment>
<ID>143</ID>
<points>-909.5,-4910.5,-726.5,-4910.5</points>
<connection>
<GID>2464</GID>
<name>clear</name></connection>
<intersection>-909.5 154</intersection>
<intersection>-900.5 155</intersection>
<intersection>-892 156</intersection>
<intersection>-884.5 157</intersection>
<intersection>-871.5 158</intersection>
<intersection>-726.5 139</intersection></hsegment>
<vsegment>
<ID>154</ID>
<points>-909.5,-4910.5,-909.5,-4865.5</points>
<connection>
<GID>2470</GID>
<name>clear</name></connection>
<intersection>-4910.5 143</intersection></vsegment>
<vsegment>
<ID>155</ID>
<points>-900.5,-4910.5,-900.5,-4873</points>
<connection>
<GID>2469</GID>
<name>clear</name></connection>
<intersection>-4910.5 143</intersection></vsegment>
<vsegment>
<ID>156</ID>
<points>-892,-4910.5,-892,-4880.5</points>
<connection>
<GID>2468</GID>
<name>clear</name></connection>
<intersection>-4910.5 143</intersection></vsegment>
<vsegment>
<ID>157</ID>
<points>-884.5,-4910.5,-884.5,-4889.5</points>
<connection>
<GID>2466</GID>
<name>clear</name></connection>
<intersection>-4910.5 143</intersection></vsegment>
<vsegment>
<ID>158</ID>
<points>-871.5,-4910.5,-871.5,-4900.5</points>
<connection>
<GID>2465</GID>
<name>clear</name></connection>
<intersection>-4910.5 143</intersection></vsegment></shape></wire>
<wire>
<ID>2654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-783,-3647,-783,-3646.5</points>
<intersection>-3647 1</intersection>
<intersection>-3646.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-787.5,-3647,-783,-3647</points>
<connection>
<GID>1861</GID>
<name>OUT</name></connection>
<intersection>-783 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-783,-3646.5,-778.5,-3646.5</points>
<connection>
<GID>1913</GID>
<name>IN_0</name></connection>
<intersection>-783 0</intersection></hsegment></shape></wire>
<wire>
<ID>2655</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-827,-3652.5,-658.5,-3652.5</points>
<intersection>-827 12</intersection>
<intersection>-802 5</intersection>
<intersection>-778.5 2</intersection>
<intersection>-658.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-778.5,-3652.5,-778.5,-3648.5</points>
<connection>
<GID>1913</GID>
<name>IN_1</name></connection>
<intersection>-3652.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-658.5,-3652.5,-658.5,-3635.5</points>
<connection>
<GID>1916</GID>
<name>IN_1</name></connection>
<intersection>-3652.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-802,-3655,-802,-3652.5</points>
<connection>
<GID>2369</GID>
<name>J</name></connection>
<intersection>-3652.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-827,-3652.5,-827,-3650.5</points>
<connection>
<GID>2296</GID>
<name>OUT</name></connection>
<intersection>-3652.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-660.5,-3644,-660.5,-3635.5</points>
<connection>
<GID>1916</GID>
<name>IN_0</name></connection>
<intersection>-3644 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-772.5,-3644,-660.5,-3644</points>
<intersection>-772.5 7</intersection>
<intersection>-763.5 2</intersection>
<intersection>-660.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-763.5,-3647,-763.5,-3644</points>
<connection>
<GID>1946</GID>
<name>N_in0</name></connection>
<intersection>-3644 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-772.5,-3647.5,-772.5,-3644</points>
<connection>
<GID>1913</GID>
<name>OUT</name></connection>
<intersection>-3644 1</intersection></vsegment></shape></wire>
<wire>
<ID>2657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1085.5,-3274.5,-1085.5,-3261.5</points>
<intersection>-3274.5 1</intersection>
<intersection>-3261.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1088.5,-3274.5,-1085.5,-3274.5</points>
<connection>
<GID>2257</GID>
<name>K</name></connection>
<intersection>-1085.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1095,-3261.5,-1085.5,-3261.5</points>
<connection>
<GID>2269</GID>
<name>OUT_0</name></connection>
<intersection>-1085.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-886,-4984,-851.5,-4984</points>
<connection>
<GID>1981</GID>
<name>IN_1</name></connection>
<intersection>-851.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-851.5,-4984,-851.5,-4983</points>
<connection>
<GID>1988</GID>
<name>OUT</name></connection>
<intersection>-4984 1</intersection></vsegment></shape></wire>
<wire>
<ID>2659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-833.5,-4973,-833.5,-4956</points>
<connection>
<GID>2478</GID>
<name>clear</name></connection>
<intersection>-4973 1</intersection>
<intersection>-4956.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-875.5,-4973,-833.5,-4973</points>
<connection>
<GID>1979</GID>
<name>Q</name></connection>
<intersection>-833.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-833.5,-4956.5,-765.5,-4956.5</points>
<connection>
<GID>2445</GID>
<name>clear</name></connection>
<connection>
<GID>2444</GID>
<name>clear</name></connection>
<connection>
<GID>2443</GID>
<name>clear</name></connection>
<connection>
<GID>2442</GID>
<name>clear</name></connection>
<connection>
<GID>2441</GID>
<name>clear</name></connection>
<intersection>-833.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-819,-4713.5,-819,-4688.5</points>
<connection>
<GID>2419</GID>
<name>IN_0</name></connection>
<intersection>-4688.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-819,-4688.5,-766.5,-4688.5</points>
<connection>
<GID>2040</GID>
<name>OUT</name></connection>
<intersection>-819 0</intersection></hsegment></shape></wire>
<wire>
<ID>2661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-866,-3616.5,-866,-3605</points>
<connection>
<GID>2196</GID>
<name>clear</name></connection>
<intersection>-3616.5 7</intersection>
<intersection>-3605.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-866,-3605.5,-798,-3605.5</points>
<connection>
<GID>2249</GID>
<name>clear</name></connection>
<connection>
<GID>2242</GID>
<name>clear</name></connection>
<connection>
<GID>2237</GID>
<name>clear</name></connection>
<connection>
<GID>2230</GID>
<name>clear</name></connection>
<connection>
<GID>2221</GID>
<name>clear</name></connection>
<intersection>-866 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-888.5,-3616.5,-866,-3616.5</points>
<connection>
<GID>2035</GID>
<name>Q</name></connection>
<intersection>-866 0</intersection></hsegment></shape></wire>
<wire>
<ID>2662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1362,-3192.5,-1362,-3192</points>
<intersection>-3192.5 2</intersection>
<intersection>-3192 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1362,-3192,-1357.5,-3192</points>
<connection>
<GID>2032</GID>
<name>IN_1</name></connection>
<intersection>-1362 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1367,-3192.5,-1362,-3192.5</points>
<connection>
<GID>2286</GID>
<name>OUT_0</name></connection>
<intersection>-1362 0</intersection></hsegment></shape></wire>
<wire>
<ID>2663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-957.5,-3635,-957.5,-3626.5</points>
<intersection>-3635 1</intersection>
<intersection>-3626.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-957.5,-3635,-955,-3635</points>
<connection>
<GID>2037</GID>
<name>OUT</name></connection>
<intersection>-957.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-957.5,-3626.5,-909.5,-3626.5</points>
<connection>
<GID>2041</GID>
<name>IN_0</name></connection>
<intersection>-957.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2664</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-909.5,-3622.5,-891.5,-3622.5</points>
<connection>
<GID>2041</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2035</GID>
<name>clear</name></connection>
<intersection>-909.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-909.5,-3622.5,-909.5,-3616.5</points>
<intersection>-3622.5 1</intersection>
<intersection>-3616.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-909.5,-3616.5,-894.5,-3616.5</points>
<connection>
<GID>2035</GID>
<name>J</name></connection>
<intersection>-909.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2665</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-888.5,-3620.5,-885.5,-3620.5</points>
<connection>
<GID>2035</GID>
<name>nQ</name></connection>
<connection>
<GID>2043</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1351,-3202,-1351,-3191</points>
<intersection>-3202 1</intersection>
<intersection>-3191 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1361.5,-3202,-1351,-3202</points>
<intersection>-1361.5 3</intersection>
<intersection>-1351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1351.5,-3191,-1351,-3191</points>
<connection>
<GID>2032</GID>
<name>OUT</name></connection>
<intersection>-1351 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1361.5,-3204.5,-1361.5,-3202</points>
<connection>
<GID>2328</GID>
<name>IN_0</name></connection>
<intersection>-3202 1</intersection></vsegment></shape></wire>
<wire>
<ID>2667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-917.5,-3661,-917.5,-3477</points>
<connection>
<GID>2045</GID>
<name>OUT_0</name></connection>
<intersection>-3661 2</intersection>
<intersection>-3630 1</intersection>
<intersection>-3629 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-938,-3630,-917.5,-3630</points>
<connection>
<GID>2047</GID>
<name>IN_1</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-917.5,-3661,-799,-3661</points>
<connection>
<GID>2369</GID>
<name>clear</name></connection>
<intersection>-917.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-917.5,-3629,-448,-3629</points>
<intersection>-917.5 0</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-448,-4980.5,-448,-3629</points>
<intersection>-4980.5 5</intersection>
<intersection>-4788.5 6</intersection>
<intersection>-4554 11</intersection>
<intersection>-4329 15</intersection>
<intersection>-4132.5 18</intersection>
<intersection>-3947 21</intersection>
<intersection>-3778 24</intersection>
<intersection>-3629 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-845.5,-4980.5,-448,-4980.5</points>
<intersection>-845.5 10</intersection>
<intersection>-448 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-864.5,-4788.5,-448,-4788.5</points>
<connection>
<GID>2056</GID>
<name>clear</name></connection>
<intersection>-864.5 7</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-864.5,-4788.5,-864.5,-4753.5</points>
<intersection>-4788.5 6</intersection>
<intersection>-4753.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-868,-4753.5,-864.5,-4753.5</points>
<connection>
<GID>1977</GID>
<name>IN_1</name></connection>
<intersection>-864.5 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-845.5,-4982,-845.5,-4980.5</points>
<connection>
<GID>1988</GID>
<name>IN_1</name></connection>
<intersection>-4980.5 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-866.5,-4554,-448,-4554</points>
<connection>
<GID>2033</GID>
<name>clear</name></connection>
<intersection>-866.5 12</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-866.5,-4554,-866.5,-4520</points>
<intersection>-4554 11</intersection>
<intersection>-4520 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-870,-4520,-866.5,-4520</points>
<connection>
<GID>1960</GID>
<name>IN_1</name></connection>
<intersection>-866.5 12</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-865.5,-4329,-448,-4329</points>
<connection>
<GID>1989</GID>
<name>clear</name></connection>
<intersection>-865.5 16</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-865.5,-4329,-865.5,-4297</points>
<intersection>-4329 15</intersection>
<intersection>-4297 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-868.5,-4297,-865.5,-4297</points>
<connection>
<GID>1901</GID>
<name>IN_1</name></connection>
<intersection>-865.5 16</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-883,-4132.5,-448,-4132.5</points>
<connection>
<GID>1965</GID>
<name>clear</name></connection>
<intersection>-883 19</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-883,-4132.5,-883,-4088.5</points>
<intersection>-4132.5 18</intersection>
<intersection>-4088.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-886.5,-4088.5,-883,-4088.5</points>
<connection>
<GID>1888</GID>
<name>IN_1</name></connection>
<intersection>-883 19</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-882,-3947,-448,-3947</points>
<connection>
<GID>1904</GID>
<name>clear</name></connection>
<intersection>-882 22</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-882,-3947,-882,-3921</points>
<intersection>-3947 21</intersection>
<intersection>-3921 23</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>-885.5,-3921,-882,-3921</points>
<connection>
<GID>2065</GID>
<name>IN_1</name></connection>
<intersection>-882 22</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-902.5,-3778,-448,-3778</points>
<connection>
<GID>1864</GID>
<name>clear</name></connection>
<intersection>-902.5 25</intersection>
<intersection>-448 4</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-902.5,-3778,-902.5,-3752</points>
<intersection>-3778 24</intersection>
<intersection>-3752 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-949.5,-3752,-902.5,-3752</points>
<connection>
<GID>2054</GID>
<name>IN_1</name></connection>
<intersection>-902.5 25</intersection></hsegment></shape></wire>
<wire>
<ID>2668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-949,-3634,-946.5,-3634</points>
<connection>
<GID>2037</GID>
<name>IN_1</name></connection>
<intersection>-946.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-946.5,-3634,-946.5,-3631</points>
<intersection>-3634 1</intersection>
<intersection>-3631 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-946.5,-3631,-944,-3631</points>
<connection>
<GID>2047</GID>
<name>OUT</name></connection>
<intersection>-946.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-971.5,-3754,-967.5,-3754</points>
<connection>
<GID>2050</GID>
<name>IN_0</name></connection>
<connection>
<GID>2049</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2670</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-971.5,-3747,-894.5,-3747</points>
<connection>
<GID>2048</GID>
<name>clear</name></connection>
<intersection>-971.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-971.5,-3750,-971.5,-3741</points>
<connection>
<GID>2050</GID>
<name>OUT_0</name></connection>
<intersection>-3747 1</intersection>
<intersection>-3741 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-971.5,-3741,-897.5,-3741</points>
<connection>
<GID>2048</GID>
<name>J</name></connection>
<intersection>-971.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2671</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-891.5,-3745,-888.5,-3745</points>
<connection>
<GID>2048</GID>
<name>nQ</name></connection>
<connection>
<GID>2052</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2672</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-961.5,-3753,-955.5,-3753</points>
<connection>
<GID>2049</GID>
<name>IN_1</name></connection>
<connection>
<GID>2054</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-866.5,-3741,-866.5,-3730</points>
<connection>
<GID>2168</GID>
<name>clear</name></connection>
<intersection>-3741 1</intersection>
<intersection>-3730.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-891.5,-3741,-866.5,-3741</points>
<connection>
<GID>2048</GID>
<name>Q</name></connection>
<intersection>-866.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-866.5,-3730.5,-798.5,-3730.5</points>
<connection>
<GID>1921</GID>
<name>clear</name></connection>
<connection>
<GID>1920</GID>
<name>clear</name></connection>
<connection>
<GID>1919</GID>
<name>clear</name></connection>
<connection>
<GID>1917</GID>
<name>clear</name></connection>
<connection>
<GID>1915</GID>
<name>clear</name></connection>
<intersection>-866.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-936.5,-3924,-936.5,-3922</points>
<connection>
<GID>2061</GID>
<name>IN_0</name></connection>
<intersection>-3924 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-936.5,-3924,-932,-3924</points>
<connection>
<GID>2060</GID>
<name>OUT</name></connection>
<intersection>-936.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2675</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-936.5,-3918,-918.5,-3918</points>
<connection>
<GID>2061</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2058</GID>
<name>clear</name></connection>
<intersection>-936.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-936.5,-3918,-936.5,-3912</points>
<intersection>-3918 1</intersection>
<intersection>-3912 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-936.5,-3912,-921.5,-3912</points>
<connection>
<GID>2058</GID>
<name>J</name></connection>
<intersection>-936.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2676</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-915.5,-3916,-912.5,-3916</points>
<connection>
<GID>2058</GID>
<name>nQ</name></connection>
<connection>
<GID>2063</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2677</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-926,-3923,-891.5,-3923</points>
<connection>
<GID>2060</GID>
<name>IN_1</name></connection>
<intersection>-891.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-891.5,-3923,-891.5,-3922</points>
<connection>
<GID>2065</GID>
<name>OUT</name></connection>
<intersection>-3923 1</intersection></vsegment></shape></wire>
<wire>
<ID>2678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-856.5,-3912,-856.5,-3892</points>
<connection>
<GID>1956</GID>
<name>clear</name></connection>
<intersection>-3912 1</intersection>
<intersection>-3892.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-915.5,-3912,-856.5,-3912</points>
<connection>
<GID>2058</GID>
<name>Q</name></connection>
<intersection>-856.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-856.5,-3892.5,-788.5,-3892.5</points>
<connection>
<GID>1885</GID>
<name>clear</name></connection>
<connection>
<GID>1884</GID>
<name>clear</name></connection>
<connection>
<GID>1881</GID>
<name>clear</name></connection>
<connection>
<GID>1870</GID>
<name>clear</name></connection>
<connection>
<GID>1860</GID>
<name>clear</name></connection>
<intersection>-856.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776,-3711,-776,-3661.5</points>
<intersection>-3711 1</intersection>
<intersection>-3679 3</intersection>
<intersection>-3661.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-779,-3711,-776,-3711</points>
<connection>
<GID>2376</GID>
<name>IN_1</name></connection>
<intersection>-776 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-778,-3661.5,-776,-3661.5</points>
<connection>
<GID>2373</GID>
<name>OUT</name></connection>
<intersection>-776 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-776,-3679,-752.5,-3679</points>
<intersection>-776 0</intersection>
<intersection>-764.5 12</intersection>
<intersection>-752.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-752.5,-3708,-752.5,-3679</points>
<intersection>-3708 7</intersection>
<intersection>-3700.5 6</intersection>
<intersection>-3692.5 9</intersection>
<intersection>-3686.5 11</intersection>
<intersection>-3679 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-766,-3700.5,-752.5,-3700.5</points>
<connection>
<GID>2381</GID>
<name>IN_1</name></connection>
<intersection>-752.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-765.5,-3708,-752.5,-3708</points>
<connection>
<GID>2378</GID>
<name>IN_1</name></connection>
<intersection>-752.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-765,-3692.5,-752.5,-3692.5</points>
<connection>
<GID>2383</GID>
<name>IN_1</name></connection>
<intersection>-752.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-765,-3686.5,-752.5,-3686.5</points>
<connection>
<GID>2385</GID>
<name>IN_1</name></connection>
<intersection>-752.5 4</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-764.5,-3681,-764.5,-3679</points>
<connection>
<GID>2388</GID>
<name>IN_1</name></connection>
<intersection>-3679 3</intersection></vsegment></shape></wire>
<wire>
<ID>2680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-869.5,-3714.5,-869.5,-3712</points>
<connection>
<GID>2162</GID>
<name>IN_0</name></connection>
<intersection>-3712 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-869.5,-3712,-785,-3712</points>
<connection>
<GID>2376</GID>
<name>OUT</name></connection>
<intersection>-869.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-856,-3714.5,-856,-3709</points>
<connection>
<GID>2163</GID>
<name>IN_0</name></connection>
<intersection>-3709 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-856,-3709,-771.5,-3709</points>
<connection>
<GID>2378</GID>
<name>OUT</name></connection>
<intersection>-856 0</intersection></hsegment></shape></wire>
<wire>
<ID>2682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-843,-3714.5,-843,-3701.5</points>
<connection>
<GID>2164</GID>
<name>IN_0</name></connection>
<intersection>-3701.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-843,-3701.5,-772,-3701.5</points>
<connection>
<GID>2381</GID>
<name>OUT</name></connection>
<intersection>-843 0</intersection></hsegment></shape></wire>
<wire>
<ID>2683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-830,-3714.5,-830,-3693.5</points>
<connection>
<GID>2165</GID>
<name>IN_0</name></connection>
<intersection>-3693.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-830,-3693.5,-771,-3693.5</points>
<connection>
<GID>2383</GID>
<name>OUT</name></connection>
<intersection>-830 0</intersection></hsegment></shape></wire>
<wire>
<ID>2684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-817.5,-3715,-817.5,-3687.5</points>
<connection>
<GID>2166</GID>
<name>IN_0</name></connection>
<intersection>-3687.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-817.5,-3687.5,-771,-3687.5</points>
<connection>
<GID>2385</GID>
<name>OUT</name></connection>
<intersection>-817.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805,-3715,-805,-3682</points>
<connection>
<GID>2167</GID>
<name>IN_0</name></connection>
<intersection>-3682 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-805,-3682,-770.5,-3682</points>
<connection>
<GID>2388</GID>
<name>OUT</name></connection>
<intersection>-805 0</intersection></hsegment></shape></wire>
<wire>
<ID>2686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-766,-3764.5,-766,-3764</points>
<intersection>-3764.5 2</intersection>
<intersection>-3764 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-768.5,-3764,-766,-3764</points>
<connection>
<GID>1867</GID>
<name>OUT</name></connection>
<intersection>-766 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-766,-3764.5,-763,-3764.5</points>
<connection>
<GID>2390</GID>
<name>IN_0</name></connection>
<intersection>-766 0</intersection></hsegment></shape></wire>
<wire>
<ID>2687</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-826,-3770.5,-644.5,-3770.5</points>
<connection>
<GID>2161</GID>
<name>OUT</name></connection>
<intersection>-811.5 6</intersection>
<intersection>-763 5</intersection>
<intersection>-644.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-644.5,-3770.5,-644.5,-3635.5</points>
<connection>
<GID>2393</GID>
<name>IN_1</name></connection>
<intersection>-3770.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-763,-3770.5,-763,-3766.5</points>
<connection>
<GID>2390</GID>
<name>IN_1</name></connection>
<intersection>-3770.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-811.5,-3772,-811.5,-3770.5</points>
<connection>
<GID>1864</GID>
<name>J</name></connection>
<intersection>-3770.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-753,-3765.5,-753,-3764</points>
<intersection>-3765.5 2</intersection>
<intersection>-3764 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-753,-3764,-646.5,-3764</points>
<connection>
<GID>1869</GID>
<name>N_in0</name></connection>
<intersection>-753 0</intersection>
<intersection>-646.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-757,-3765.5,-753,-3765.5</points>
<connection>
<GID>2390</GID>
<name>OUT</name></connection>
<intersection>-753 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-646.5,-3764,-646.5,-3635.5</points>
<connection>
<GID>2393</GID>
<name>IN_0</name></connection>
<intersection>-3764 1</intersection></vsegment></shape></wire>
<wire>
<ID>2689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-991,-3497,-991,-3496.5</points>
<connection>
<GID>2071</GID>
<name>IN_1</name></connection>
<intersection>-3496.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-994.5,-3496.5,-994.5,-3492.5</points>
<connection>
<GID>1908</GID>
<name>OUT_0</name></connection>
<intersection>-3496.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-994.5,-3496.5,-991,-3496.5</points>
<intersection>-994.5 1</intersection>
<intersection>-991 0</intersection></hsegment></shape></wire>
<wire>
<ID>2690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-989,-3497,-989,-3496.5</points>
<connection>
<GID>2071</GID>
<name>IN_0</name></connection>
<intersection>-3496.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-982.5,-3496.5,-982.5,-3492</points>
<connection>
<GID>2066</GID>
<name>OUT_0</name></connection>
<intersection>-3496.5 2</intersection>
<intersection>-3492 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-989,-3496.5,-982.5,-3496.5</points>
<intersection>-989 0</intersection>
<intersection>-982.5 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-982.5,-3492,-960.5,-3492</points>
<intersection>-982.5 1</intersection>
<intersection>-960.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-960.5,-3492,-960.5,-3490</points>
<connection>
<GID>2139</GID>
<name>N_in0</name></connection>
<intersection>-3492 4</intersection></vsegment></shape></wire>
<wire>
<ID>2691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-990,-3649,-990,-3645.5</points>
<connection>
<GID>2344</GID>
<name>OUT_0</name></connection>
<intersection>-3649 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-990,-3649,-986,-3649</points>
<connection>
<GID>2074</GID>
<name>IN_1</name></connection>
<intersection>-990 0</intersection></hsegment></shape></wire>
<wire>
<ID>2692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-984,-3649,-984,-3647</points>
<connection>
<GID>2074</GID>
<name>IN_0</name></connection>
<intersection>-3647 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-983.5,-3647,-983.5,-3645.5</points>
<connection>
<GID>2077</GID>
<name>OUT_0</name></connection>
<intersection>-3647 2</intersection>
<intersection>-3646.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-984,-3647,-983.5,-3647</points>
<intersection>-984 0</intersection>
<intersection>-983.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-983.5,-3646.5,-972.5,-3646.5</points>
<intersection>-983.5 1</intersection>
<intersection>-972.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-972.5,-3646.5,-972.5,-3644.5</points>
<connection>
<GID>2142</GID>
<name>N_in0</name></connection>
<intersection>-3646.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>2693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-999,-3772.5,-999,-3769</points>
<connection>
<GID>2088</GID>
<name>OUT_0</name></connection>
<intersection>-3772.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-999,-3772.5,-995,-3772.5</points>
<connection>
<GID>2082</GID>
<name>IN_1</name></connection>
<intersection>-999 0</intersection></hsegment></shape></wire>
<wire>
<ID>2694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-993,-3772.5,-993,-3770.5</points>
<connection>
<GID>2082</GID>
<name>IN_0</name></connection>
<intersection>-3770.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-992.5,-3770.5,-992.5,-3769</points>
<connection>
<GID>2084</GID>
<name>OUT_0</name></connection>
<intersection>-3770.5 2</intersection>
<intersection>-3769.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-993,-3770.5,-992.5,-3770.5</points>
<intersection>-993 0</intersection>
<intersection>-992.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-992.5,-3769.5,-982,-3769.5</points>
<intersection>-992.5 1</intersection>
<intersection>-982 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-982,-3769.5,-982,-3767.5</points>
<connection>
<GID>2144</GID>
<name>N_in0</name></connection>
<intersection>-3769.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>2695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-984.5,-3948.5,-984.5,-3945</points>
<connection>
<GID>2101</GID>
<name>OUT_0</name></connection>
<intersection>-3948.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-984.5,-3948.5,-981.5,-3948.5</points>
<intersection>-984.5 0</intersection>
<intersection>-981.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-981.5,-3949,-981.5,-3948.5</points>
<connection>
<GID>2089</GID>
<name>IN_1</name></connection>
<intersection>-3948.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>2696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-979.5,-3949,-979.5,-3946.5</points>
<connection>
<GID>2089</GID>
<name>IN_0</name></connection>
<intersection>-3946.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-977.5,-3946.5,-977.5,-3945</points>
<connection>
<GID>2093</GID>
<name>OUT_0</name></connection>
<intersection>-3946.5 2</intersection>
<intersection>-3945 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-979.5,-3946.5,-977.5,-3946.5</points>
<intersection>-979.5 0</intersection>
<intersection>-977.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-977.5,-3945,-966,-3945</points>
<connection>
<GID>2146</GID>
<name>N_in0</name></connection>
<intersection>-977.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-966,-4146,-966,-4142.5</points>
<connection>
<GID>2113</GID>
<name>OUT_0</name></connection>
<intersection>-4146 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-966,-4146,-962,-4146</points>
<connection>
<GID>2105</GID>
<name>IN_1</name></connection>
<intersection>-966 0</intersection></hsegment></shape></wire>
<wire>
<ID>2698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-960,-4146,-960,-4144</points>
<connection>
<GID>2105</GID>
<name>IN_0</name></connection>
<intersection>-4144 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-959.5,-4144,-959.5,-4142.5</points>
<connection>
<GID>2109</GID>
<name>OUT_0</name></connection>
<intersection>-4144 2</intersection>
<intersection>-4143 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-960,-4144,-959.5,-4144</points>
<intersection>-960 0</intersection>
<intersection>-959.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-959.5,-4143,-949,-4143</points>
<connection>
<GID>2148</GID>
<name>N_in0</name></connection>
<intersection>-959.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-972.5,-4363.5,-972.5,-4360</points>
<connection>
<GID>2121</GID>
<name>OUT_0</name></connection>
<intersection>-4363.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-972.5,-4363.5,-968.5,-4363.5</points>
<connection>
<GID>2115</GID>
<name>IN_1</name></connection>
<intersection>-972.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-966.5,-4363.5,-966.5,-4361.5</points>
<connection>
<GID>2115</GID>
<name>IN_0</name></connection>
<intersection>-4361.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-966,-4361.5,-966,-4360</points>
<connection>
<GID>2117</GID>
<name>OUT_0</name></connection>
<intersection>-4361.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-966.5,-4361.5,-956.5,-4361.5</points>
<connection>
<GID>2150</GID>
<name>N_in0</name></connection>
<intersection>-966.5 0</intersection>
<intersection>-966 1</intersection></hsegment></shape></wire>
<wire>
<ID>2701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-971.5,-4605.5,-971.5,-4602</points>
<connection>
<GID>2128</GID>
<name>OUT_0</name></connection>
<intersection>-4605.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-971.5,-4605.5,-967.5,-4605.5</points>
<connection>
<GID>2122</GID>
<name>IN_1</name></connection>
<intersection>-971.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-965.5,-4605.5,-965.5,-4603.5</points>
<connection>
<GID>2122</GID>
<name>IN_0</name></connection>
<intersection>-4603.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-965,-4603.5,-965,-4602</points>
<connection>
<GID>2124</GID>
<name>OUT_0</name></connection>
<intersection>-4603.5 2</intersection>
<intersection>-4602.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-965.5,-4603.5,-965,-4603.5</points>
<intersection>-965.5 0</intersection>
<intersection>-965 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-965,-4602.5,-955,-4602.5</points>
<connection>
<GID>2152</GID>
<name>N_in0</name></connection>
<intersection>-965 1</intersection></hsegment></shape></wire>
<wire>
<ID>2703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-964.5,-4819,-964.5,-4815.5</points>
<connection>
<GID>2136</GID>
<name>OUT_0</name></connection>
<intersection>-4819 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-964.5,-4819,-960.5,-4819</points>
<connection>
<GID>2130</GID>
<name>IN_1</name></connection>
<intersection>-964.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-958.5,-4819,-958.5,-4817</points>
<connection>
<GID>2130</GID>
<name>IN_0</name></connection>
<intersection>-4817 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-958,-4817,-958,-4815.5</points>
<connection>
<GID>2132</GID>
<name>OUT_0</name></connection>
<intersection>-4817 2</intersection>
<intersection>-4816.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-958.5,-4817,-958,-4817</points>
<intersection>-958.5 0</intersection>
<intersection>-958 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-958,-4816.5,-949,-4816.5</points>
<connection>
<GID>2154</GID>
<name>N_in0</name></connection>
<intersection>-958 1</intersection></hsegment></shape></wire>
<wire>
<ID>2156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-802,-3646,-802,-3634</points>
<intersection>-3646 1</intersection>
<intersection>-3634 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-802,-3646,-793.5,-3646</points>
<connection>
<GID>1861</GID>
<name>IN_0</name></connection>
<intersection>-802 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-810.5,-3634,-802,-3634</points>
<intersection>-810.5 15</intersection>
<intersection>-802 0</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-810.5,-3640.5,-810.5,-3634</points>
<connection>
<GID>1961</GID>
<name>OUT</name></connection>
<intersection>-3634 2</intersection></vsegment></shape></wire>
<wire>
<ID>2157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-798.5,-3778,-798.5,-3772</points>
<intersection>-3778 2</intersection>
<intersection>-3772 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-805.5,-3772,-798.5,-3772</points>
<connection>
<GID>1864</GID>
<name>Q</name></connection>
<intersection>-798.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-798.5,-3778,-791.5,-3778</points>
<connection>
<GID>1868</GID>
<name>IN_0</name></connection>
<intersection>-798.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-797,-3930,-797,-3927.5</points>
<intersection>-3930 2</intersection>
<intersection>-3927.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-801,-3927.5,-797,-3927.5</points>
<connection>
<GID>1943</GID>
<name>OUT</name></connection>
<intersection>-797 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-797,-3930,-792.5,-3930</points>
<connection>
<GID>1863</GID>
<name>IN_0</name></connection>
<intersection>-797 0</intersection></hsegment></shape></wire>
<wire>
<ID>2159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-659.5,-3629.5,-659.5,-3624.5</points>
<connection>
<GID>1916</GID>
<name>OUT</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-643.5,-3624.5,-643.5,-3619.5</points>
<connection>
<GID>1866</GID>
<name>IN_0</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-659.5,-3624.5,-643.5,-3624.5</points>
<intersection>-659.5 0</intersection>
<intersection>-643.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-778.5,-3763,-778.5,-3757.5</points>
<intersection>-3763 2</intersection>
<intersection>-3757.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-782.5,-3757.5,-778.5,-3757.5</points>
<connection>
<GID>1865</GID>
<name>OUT</name></connection>
<intersection>-778.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-778.5,-3763,-774.5,-3763</points>
<connection>
<GID>1867</GID>
<name>IN_0</name></connection>
<intersection>-778.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776.5,-3860,-776.5,-3779</points>
<intersection>-3860 2</intersection>
<intersection>-3805.5 3</intersection>
<intersection>-3779 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-785.5,-3779,-776.5,-3779</points>
<connection>
<GID>1868</GID>
<name>OUT</name></connection>
<intersection>-776.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-777.5,-3860,-776.5,-3860</points>
<connection>
<GID>1873</GID>
<name>IN_1</name></connection>
<intersection>-776.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-776.5,-3805.5,-756,-3805.5</points>
<intersection>-776.5 0</intersection>
<intersection>-756 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-756,-3854.5,-756,-3805.5</points>
<intersection>-3854.5 5</intersection>
<intersection>-3846.5 6</intersection>
<intersection>-3838.5 7</intersection>
<intersection>-3828 8</intersection>
<intersection>-3817 9</intersection>
<intersection>-3805.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-762,-3854.5,-756,-3854.5</points>
<connection>
<GID>1877</GID>
<name>IN_1</name></connection>
<intersection>-756 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-761.5,-3846.5,-756,-3846.5</points>
<connection>
<GID>1882</GID>
<name>IN_1</name></connection>
<intersection>-756 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-760.5,-3838.5,-756,-3838.5</points>
<connection>
<GID>1887</GID>
<name>IN_1</name></connection>
<intersection>-756 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-760,-3828,-756,-3828</points>
<connection>
<GID>1889</GID>
<name>IN_1</name></connection>
<intersection>-756 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-760.5,-3817,-756,-3817</points>
<connection>
<GID>1894</GID>
<name>IN_1</name></connection>
<intersection>-756 4</intersection></hsegment></shape></wire>
<wire>
<ID>2162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-793,-4109.5,-786,-4109.5</points>
<connection>
<GID>2020</GID>
<name>OUT</name></connection>
<connection>
<GID>1874</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-645.5,-3629.5,-645.5,-3624.5</points>
<connection>
<GID>2393</GID>
<name>OUT</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-641.5,-3624.5,-641.5,-3619.5</points>
<connection>
<GID>1866</GID>
<name>IN_1</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-645.5,-3624.5,-641.5,-3624.5</points>
<intersection>-645.5 0</intersection>
<intersection>-641.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-782.5,-4308.5,-778,-4308.5</points>
<connection>
<GID>2133</GID>
<name>OUT</name></connection>
<connection>
<GID>1876</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-937.5,-4091.5,-937.5,-4089.5</points>
<connection>
<GID>1875</GID>
<name>IN_0</name></connection>
<intersection>-4091.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-937.5,-4091.5,-933,-4091.5</points>
<connection>
<GID>1872</GID>
<name>OUT</name></connection>
<intersection>-937.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-789,-4530.5,-782.5,-4530.5</points>
<connection>
<GID>2382</GID>
<name>OUT</name></connection>
<connection>
<GID>1880</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-937.5,-4085.5,-919.5,-4085.5</points>
<connection>
<GID>1875</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1871</GID>
<name>clear</name></connection>
<intersection>-937.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-937.5,-4085.5,-937.5,-4079.5</points>
<intersection>-4085.5 1</intersection>
<intersection>-4079.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-937.5,-4079.5,-922.5,-4079.5</points>
<connection>
<GID>1871</GID>
<name>J</name></connection>
<intersection>-937.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-787,-4764.5,-781,-4764.5</points>
<connection>
<GID>2429</GID>
<name>OUT</name></connection>
<connection>
<GID>1883</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2169</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-916.5,-4083.5,-913.5,-4083.5</points>
<connection>
<GID>1871</GID>
<name>nQ</name></connection>
<connection>
<GID>1879</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-778,-4991.5,-772,-4991.5</points>
<connection>
<GID>2467</GID>
<name>OUT</name></connection>
<connection>
<GID>1893</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-859.5,-3876.5,-859.5,-3861</points>
<connection>
<GID>1930</GID>
<name>IN_0</name></connection>
<intersection>-3861 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-859.5,-3861,-783.5,-3861</points>
<connection>
<GID>1873</GID>
<name>OUT</name></connection>
<intersection>-859.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-846,-3876.5,-846,-3855.5</points>
<connection>
<GID>1931</GID>
<name>IN_0</name></connection>
<intersection>-3855.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-846,-3855.5,-768,-3855.5</points>
<connection>
<GID>1877</GID>
<name>OUT</name></connection>
<intersection>-846 0</intersection></hsegment></shape></wire>
<wire>
<ID>2173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-833,-3876.5,-833,-3847.5</points>
<connection>
<GID>1932</GID>
<name>IN_0</name></connection>
<intersection>-3847.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-833,-3847.5,-767.5,-3847.5</points>
<connection>
<GID>1882</GID>
<name>OUT</name></connection>
<intersection>-833 0</intersection></hsegment></shape></wire>
<wire>
<ID>2174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-980.5,-3932,-980.5,-3778.5</points>
<intersection>-3932 13</intersection>
<intersection>-3839.5 1</intersection>
<intersection>-3829.5 3</intersection>
<intersection>-3818.5 5</intersection>
<intersection>-3809.5 7</intersection>
<intersection>-3802 9</intersection>
<intersection>-3794.5 11</intersection>
<intersection>-3780 15</intersection>
<intersection>-3778.5 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-980.5,-3839.5,-949.5,-3839.5</points>
<connection>
<GID>1950</GID>
<name>IN_0</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-980.5,-3829.5,-950,-3829.5</points>
<connection>
<GID>1951</GID>
<name>IN_0</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-980.5,-3818.5,-951.5,-3818.5</points>
<connection>
<GID>1952</GID>
<name>IN_0</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-980.5,-3809.5,-952,-3809.5</points>
<connection>
<GID>1953</GID>
<name>IN_0</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-980.5,-3802,-953,-3802</points>
<connection>
<GID>1954</GID>
<name>IN_0</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-980.5,-3794.5,-954,-3794.5</points>
<connection>
<GID>1955</GID>
<name>IN_0</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-980.5,-3932,-792.5,-3932</points>
<connection>
<GID>1863</GID>
<name>IN_1</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-980.5,-3780,-791.5,-3780</points>
<connection>
<GID>1868</GID>
<name>IN_1</name></connection>
<intersection>-980.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-994,-3778.5,-980.5,-3778.5</points>
<connection>
<GID>2082</GID>
<name>OUT</name></connection>
<intersection>-980.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-820,-3876.5,-820,-3839.5</points>
<connection>
<GID>1933</GID>
<name>IN_0</name></connection>
<intersection>-3839.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-820,-3839.5,-766.5,-3839.5</points>
<connection>
<GID>1887</GID>
<name>OUT</name></connection>
<intersection>-820 0</intersection></hsegment></shape></wire>
<wire>
<ID>2176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-807.5,-3877,-807.5,-3829</points>
<connection>
<GID>1934</GID>
<name>IN_0</name></connection>
<intersection>-3829 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-807.5,-3829,-766,-3829</points>
<connection>
<GID>1889</GID>
<name>OUT</name></connection>
<intersection>-807.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-790,-3660.5,-790,-3655</points>
<intersection>-3660.5 2</intersection>
<intersection>-3655 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-796,-3655,-790,-3655</points>
<connection>
<GID>2369</GID>
<name>Q</name></connection>
<intersection>-790 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-790,-3660.5,-784,-3660.5</points>
<connection>
<GID>2373</GID>
<name>IN_0</name></connection>
<intersection>-790 0</intersection></hsegment></shape></wire>
<wire>
<ID>2178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795,-3877,-795,-3818</points>
<connection>
<GID>1936</GID>
<name>IN_0</name></connection>
<intersection>-3818 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-795,-3818,-766.5,-3818</points>
<connection>
<GID>1894</GID>
<name>OUT</name></connection>
<intersection>-795 0</intersection></hsegment></shape></wire>
<wire>
<ID>2179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-625,-3937.5,-625,-3635.5</points>
<connection>
<GID>1896</GID>
<name>IN_1</name></connection>
<intersection>-3937.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-817.5,-3937.5,-625,-3937.5</points>
<connection>
<GID>1924</GID>
<name>OUT</name></connection>
<intersection>-817.5 5</intersection>
<intersection>-779.5 4</intersection>
<intersection>-625 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-779.5,-3937.5,-779.5,-3933</points>
<connection>
<GID>1900</GID>
<name>IN_1</name></connection>
<intersection>-3937.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-817.5,-3941,-817.5,-3937.5</points>
<intersection>-3941 6</intersection>
<intersection>-3937.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-817.5,-3941,-805.5,-3941</points>
<connection>
<GID>1904</GID>
<name>J</name></connection>
<intersection>-817.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>2180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-626,-3629.5,-626,-3624.5</points>
<connection>
<GID>1896</GID>
<name>OUT</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-639.5,-3624.5,-639.5,-3619.5</points>
<connection>
<GID>1866</GID>
<name>IN_2</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-639.5,-3624.5,-626,-3624.5</points>
<intersection>-639.5 1</intersection>
<intersection>-626 0</intersection></hsegment></shape></wire>
<wire>
<ID>2181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-609.5,-3630,-609.5,-3624.5</points>
<connection>
<GID>1972</GID>
<name>OUT</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-637.5,-3624.5,-637.5,-3619.5</points>
<connection>
<GID>1866</GID>
<name>IN_3</name></connection>
<intersection>-3624.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-637.5,-3624.5,-609.5,-3624.5</points>
<intersection>-637.5 1</intersection>
<intersection>-609.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-927,-4090.5,-892.5,-4090.5</points>
<connection>
<GID>1872</GID>
<name>IN_1</name></connection>
<intersection>-892.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-892.5,-4090.5,-892.5,-4089.5</points>
<connection>
<GID>1888</GID>
<name>OUT</name></connection>
<intersection>-4090.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-786.5,-3931,-779.5,-3931</points>
<connection>
<GID>1863</GID>
<name>OUT</name></connection>
<connection>
<GID>1900</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-766.5,-3926,-766.5,-3925</points>
<intersection>-3926 1</intersection>
<intersection>-3925 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-766.5,-3926,-627,-3926</points>
<connection>
<GID>1902</GID>
<name>N_in0</name></connection>
<intersection>-766.5 0</intersection>
<intersection>-627 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-772,-3925,-766.5,-3925</points>
<intersection>-772 6</intersection>
<intersection>-766.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-627,-3926,-627,-3635.5</points>
<connection>
<GID>1896</GID>
<name>IN_0</name></connection>
<intersection>-3926 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-772,-3932,-772,-3925</points>
<intersection>-3932 7</intersection>
<intersection>-3925 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-773.5,-3932,-772,-3932</points>
<connection>
<GID>1900</GID>
<name>OUT</name></connection>
<intersection>-772 6</intersection></hsegment></shape></wire>
<wire>
<ID>2185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-870.5,-3724,-870.5,-3720.5</points>
<connection>
<GID>2162</GID>
<name>OUT</name></connection>
<intersection>-3724 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-870.5,-3724,-869.5,-3724</points>
<connection>
<GID>2168</GID>
<name>IN_0</name></connection>
<intersection>-870.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-857,-3724.5,-857,-3720.5</points>
<connection>
<GID>2163</GID>
<name>OUT</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-857,-3724.5,-853.5,-3724.5</points>
<connection>
<GID>1915</GID>
<name>IN_0</name></connection>
<intersection>-857 0</intersection></hsegment></shape></wire>
<wire>
<ID>2187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844,-3724.5,-844,-3720.5</points>
<connection>
<GID>2164</GID>
<name>OUT</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-844,-3724.5,-840,-3724.5</points>
<connection>
<GID>1917</GID>
<name>IN_0</name></connection>
<intersection>-844 0</intersection></hsegment></shape></wire>
<wire>
<ID>2188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-828,-3724.5,-828,-3720.5</points>
<intersection>-3724.5 1</intersection>
<intersection>-3720.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-828,-3724.5,-825,-3724.5</points>
<connection>
<GID>1919</GID>
<name>IN_0</name></connection>
<intersection>-828 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-831,-3720.5,-828,-3720.5</points>
<connection>
<GID>2165</GID>
<name>OUT</name></connection>
<intersection>-828 0</intersection></hsegment></shape></wire>
<wire>
<ID>2189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-818.5,-3723,-818.5,-3721</points>
<connection>
<GID>2166</GID>
<name>OUT</name></connection>
<intersection>-3723 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-818.5,-3723,-814.5,-3723</points>
<intersection>-818.5 0</intersection>
<intersection>-814.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-814.5,-3724.5,-814.5,-3723</points>
<connection>
<GID>1920</GID>
<name>IN_0</name></connection>
<intersection>-3723 1</intersection></vsegment></shape></wire>
<wire>
<ID>2190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-806,-3723,-806,-3721</points>
<connection>
<GID>2167</GID>
<name>OUT</name></connection>
<intersection>-3723 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-806,-3723,-801.5,-3723</points>
<intersection>-806 0</intersection>
<intersection>-801.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-801.5,-3724.5,-801.5,-3723</points>
<connection>
<GID>1921</GID>
<name>IN_0</name></connection>
<intersection>-3723 1</intersection></vsegment></shape></wire>
<wire>
<ID>2191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-859.5,-3732,-859.5,-3724</points>
<connection>
<GID>1923</GID>
<name>IN_0</name></connection>
<intersection>-3724 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-863.5,-3724,-859.5,-3724</points>
<connection>
<GID>2168</GID>
<name>OUT_0</name></connection>
<intersection>-859.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844.5,-3732,-844.5,-3724.5</points>
<connection>
<GID>1925</GID>
<name>IN_0</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-847.5,-3724.5,-844.5,-3724.5</points>
<connection>
<GID>1915</GID>
<name>OUT_0</name></connection>
<intersection>-844.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-829.5,-3732,-829.5,-3724.5</points>
<connection>
<GID>1926</GID>
<name>IN_0</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-834,-3724.5,-829.5,-3724.5</points>
<connection>
<GID>1917</GID>
<name>OUT_0</name></connection>
<intersection>-829.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-818,-3731.5,-818,-3724.5</points>
<connection>
<GID>1927</GID>
<name>IN_0</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-819,-3724.5,-818,-3724.5</points>
<connection>
<GID>1919</GID>
<name>OUT_0</name></connection>
<intersection>-818 0</intersection></hsegment></shape></wire>
<wire>
<ID>2195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805,-3732,-805,-3724.5</points>
<connection>
<GID>1928</GID>
<name>IN_0</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-808.5,-3724.5,-805,-3724.5</points>
<connection>
<GID>1920</GID>
<name>OUT_0</name></connection>
<intersection>-805 0</intersection></hsegment></shape></wire>
<wire>
<ID>2196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-792,-3731.5,-792,-3724.5</points>
<connection>
<GID>1929</GID>
<name>IN_0</name></connection>
<intersection>-3724.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-795.5,-3724.5,-792,-3724.5</points>
<connection>
<GID>1921</GID>
<name>OUT_0</name></connection>
<intersection>-792 0</intersection></hsegment></shape></wire>
<wire>
<ID>2197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-859.5,-3741.5,-859.5,-3736</points>
<connection>
<GID>1923</GID>
<name>OUT_0</name></connection>
<intersection>-3741.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-844.5,-3747.5,-844.5,-3741.5</points>
<connection>
<GID>2159</GID>
<name>IN_3</name></connection>
<intersection>-3741.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-859.5,-3741.5,-844.5,-3741.5</points>
<intersection>-859.5 0</intersection>
<intersection>-844.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844.5,-3741,-844.5,-3736</points>
<connection>
<GID>1925</GID>
<name>OUT_0</name></connection>
<intersection>-3741 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-842.5,-3747.5,-842.5,-3741</points>
<connection>
<GID>2159</GID>
<name>IN_2</name></connection>
<intersection>-3741 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-844.5,-3741,-842.5,-3741</points>
<intersection>-844.5 0</intersection>
<intersection>-842.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-829.5,-3741.5,-829.5,-3736</points>
<connection>
<GID>1926</GID>
<name>OUT_0</name></connection>
<intersection>-3741.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-840.5,-3747.5,-840.5,-3741.5</points>
<connection>
<GID>2159</GID>
<name>IN_1</name></connection>
<intersection>-3741.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-840.5,-3741.5,-829.5,-3741.5</points>
<intersection>-840.5 1</intersection>
<intersection>-829.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-818,-3742.5,-818,-3735.5</points>
<connection>
<GID>1927</GID>
<name>OUT_0</name></connection>
<intersection>-3742.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-838.5,-3747.5,-838.5,-3742.5</points>
<connection>
<GID>2159</GID>
<name>IN_0</name></connection>
<intersection>-3742.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-838.5,-3742.5,-818,-3742.5</points>
<intersection>-838.5 1</intersection>
<intersection>-818 0</intersection></hsegment></shape></wire>
<wire>
<ID>2201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-793,-3946,-793,-3941</points>
<intersection>-3946 2</intersection>
<intersection>-3941 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-799.5,-3941,-793,-3941</points>
<connection>
<GID>1904</GID>
<name>Q</name></connection>
<intersection>-793 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-793,-3946,-786,-3946</points>
<connection>
<GID>1935</GID>
<name>IN_0</name></connection>
<intersection>-793 0</intersection></hsegment></shape></wire>
<wire>
<ID>2202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-860.5,-3886,-860.5,-3882.5</points>
<connection>
<GID>1930</GID>
<name>OUT</name></connection>
<intersection>-3886 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-860.5,-3886,-859.5,-3886</points>
<connection>
<GID>1956</GID>
<name>IN_0</name></connection>
<intersection>-860.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-851.5,-4058.5,-851.5,-4043</points>
<connection>
<GID>2008</GID>
<name>IN_0</name></connection>
<intersection>-4043 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-851.5,-4043,-781,-4043</points>
<connection>
<GID>1939</GID>
<name>OUT</name></connection>
<intersection>-851.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-774,-4042,-774,-3947</points>
<intersection>-4042 2</intersection>
<intersection>-3980 3</intersection>
<intersection>-3947 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-780,-3947,-774,-3947</points>
<connection>
<GID>1935</GID>
<name>OUT</name></connection>
<intersection>-774 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-775,-4042,-774,-4042</points>
<connection>
<GID>1939</GID>
<name>IN_1</name></connection>
<intersection>-774 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-774,-3980,-761,-3980</points>
<intersection>-774 0</intersection>
<intersection>-761 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-761,-4030,-761,-3980</points>
<intersection>-4030 6</intersection>
<intersection>-4021.5 5</intersection>
<intersection>-4014 7</intersection>
<intersection>-4005 8</intersection>
<intersection>-3997 9</intersection>
<intersection>-3980 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-765,-4021.5,-761,-4021.5</points>
<connection>
<GID>1959</GID>
<name>IN_1</name></connection>
<intersection>-761 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-765,-4030,-761,-4030</points>
<connection>
<GID>1958</GID>
<name>IN_1</name></connection>
<intersection>-761 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-764,-4014,-761,-4014</points>
<connection>
<GID>1962</GID>
<name>IN_1</name></connection>
<intersection>-761 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-763.5,-4005,-761,-4005</points>
<connection>
<GID>1964</GID>
<name>IN_1</name></connection>
<intersection>-761 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-763,-3997,-761,-3997</points>
<connection>
<GID>1966</GID>
<name>IN_1</name></connection>
<intersection>-761 4</intersection></hsegment></shape></wire>
<wire>
<ID>2205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-847,-3886.5,-847,-3882.5</points>
<connection>
<GID>1931</GID>
<name>OUT</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-847,-3886.5,-843.5,-3886.5</points>
<connection>
<GID>1860</GID>
<name>IN_0</name></connection>
<intersection>-847 0</intersection></hsegment></shape></wire>
<wire>
<ID>2206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-834,-3886.5,-834,-3882.5</points>
<connection>
<GID>1932</GID>
<name>OUT</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-834,-3886.5,-830,-3886.5</points>
<connection>
<GID>1870</GID>
<name>IN_0</name></connection>
<intersection>-834 0</intersection></hsegment></shape></wire>
<wire>
<ID>2207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-838,-4058.5,-838,-4031</points>
<connection>
<GID>2009</GID>
<name>IN_0</name></connection>
<intersection>-4031 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-838,-4031,-771,-4031</points>
<connection>
<GID>1958</GID>
<name>OUT</name></connection>
<intersection>-838 0</intersection></hsegment></shape></wire>
<wire>
<ID>2208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1105,-3264,-1105,-3261.5</points>
<intersection>-3264 2</intersection>
<intersection>-3261.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1105,-3261.5,-1101,-3261.5</points>
<connection>
<GID>2269</GID>
<name>IN_0</name></connection>
<intersection>-1105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1108.5,-3264,-1105,-3264</points>
<connection>
<GID>2310</GID>
<name>OUT</name></connection>
<intersection>-1105 0</intersection></hsegment></shape></wire>
<wire>
<ID>2209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-818,-3886.5,-818,-3882.5</points>
<intersection>-3886.5 1</intersection>
<intersection>-3882.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-818,-3886.5,-815,-3886.5</points>
<connection>
<GID>1881</GID>
<name>IN_0</name></connection>
<intersection>-818 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-821,-3882.5,-818,-3882.5</points>
<connection>
<GID>1933</GID>
<name>OUT</name></connection>
<intersection>-818 0</intersection></hsegment></shape></wire>
<wire>
<ID>2210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808.5,-3885,-808.5,-3883</points>
<connection>
<GID>1934</GID>
<name>OUT</name></connection>
<intersection>-3885 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-808.5,-3885,-804.5,-3885</points>
<intersection>-808.5 0</intersection>
<intersection>-804.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-804.5,-3886.5,-804.5,-3885</points>
<connection>
<GID>1884</GID>
<name>IN_0</name></connection>
<intersection>-3885 1</intersection></vsegment></shape></wire>
<wire>
<ID>2211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-796,-3885,-796,-3883</points>
<connection>
<GID>1936</GID>
<name>OUT</name></connection>
<intersection>-3885 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-796,-3885,-791.5,-3885</points>
<intersection>-796 0</intersection>
<intersection>-791.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-791.5,-3886.5,-791.5,-3885</points>
<connection>
<GID>1885</GID>
<name>IN_0</name></connection>
<intersection>-3885 1</intersection></vsegment></shape></wire>
<wire>
<ID>2212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-849.5,-3894,-849.5,-3886</points>
<connection>
<GID>1890</GID>
<name>IN_0</name></connection>
<intersection>-3886 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-853.5,-3886,-849.5,-3886</points>
<connection>
<GID>1956</GID>
<name>OUT_0</name></connection>
<intersection>-849.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-834.5,-3894,-834.5,-3886.5</points>
<connection>
<GID>1899</GID>
<name>IN_0</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-837.5,-3886.5,-834.5,-3886.5</points>
<connection>
<GID>1860</GID>
<name>OUT_0</name></connection>
<intersection>-834.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-819.5,-3894,-819.5,-3886.5</points>
<connection>
<GID>1905</GID>
<name>IN_0</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-824,-3886.5,-819.5,-3886.5</points>
<connection>
<GID>1870</GID>
<name>OUT_0</name></connection>
<intersection>-819.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808,-3893.5,-808,-3886.5</points>
<connection>
<GID>1907</GID>
<name>IN_0</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-809,-3886.5,-808,-3886.5</points>
<connection>
<GID>1881</GID>
<name>OUT_0</name></connection>
<intersection>-808 0</intersection></hsegment></shape></wire>
<wire>
<ID>2216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795,-3894,-795,-3886.5</points>
<connection>
<GID>1911</GID>
<name>IN_0</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-798.5,-3886.5,-795,-3886.5</points>
<connection>
<GID>1884</GID>
<name>OUT_0</name></connection>
<intersection>-795 0</intersection></hsegment></shape></wire>
<wire>
<ID>2217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-782,-3893.5,-782,-3886.5</points>
<connection>
<GID>1912</GID>
<name>IN_0</name></connection>
<intersection>-3886.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-785.5,-3886.5,-782,-3886.5</points>
<connection>
<GID>1885</GID>
<name>OUT_0</name></connection>
<intersection>-782 0</intersection></hsegment></shape></wire>
<wire>
<ID>2218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-849.5,-3903.5,-849.5,-3898</points>
<connection>
<GID>1890</GID>
<name>OUT_0</name></connection>
<intersection>-3903.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-834.5,-3909.5,-834.5,-3903.5</points>
<connection>
<GID>1914</GID>
<name>IN_3</name></connection>
<intersection>-3903.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-849.5,-3903.5,-834.5,-3903.5</points>
<intersection>-849.5 0</intersection>
<intersection>-834.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-834.5,-3903,-834.5,-3898</points>
<connection>
<GID>1899</GID>
<name>OUT_0</name></connection>
<intersection>-3903 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-832.5,-3909.5,-832.5,-3903</points>
<connection>
<GID>1914</GID>
<name>IN_2</name></connection>
<intersection>-3903 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-834.5,-3903,-832.5,-3903</points>
<intersection>-834.5 0</intersection>
<intersection>-832.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-825,-4058.5,-825,-4022.5</points>
<connection>
<GID>2010</GID>
<name>IN_0</name></connection>
<intersection>-4022.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-825,-4022.5,-771,-4022.5</points>
<connection>
<GID>1959</GID>
<name>OUT</name></connection>
<intersection>-825 0</intersection></hsegment></shape></wire>
<wire>
<ID>2221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-819.5,-3903.5,-819.5,-3898</points>
<connection>
<GID>1905</GID>
<name>OUT_0</name></connection>
<intersection>-3903.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-830.5,-3909.5,-830.5,-3903.5</points>
<connection>
<GID>1914</GID>
<name>IN_1</name></connection>
<intersection>-3903.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-830.5,-3903.5,-819.5,-3903.5</points>
<intersection>-830.5 1</intersection>
<intersection>-819.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808,-3904.5,-808,-3897.5</points>
<connection>
<GID>1907</GID>
<name>OUT_0</name></connection>
<intersection>-3904.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-828.5,-3909.5,-828.5,-3904.5</points>
<connection>
<GID>1914</GID>
<name>IN_0</name></connection>
<intersection>-3904.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-828.5,-3904.5,-808,-3904.5</points>
<intersection>-828.5 1</intersection>
<intersection>-808 0</intersection></hsegment></shape></wire>
<wire>
<ID>2223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-812,-4058.5,-812,-4015</points>
<connection>
<GID>2011</GID>
<name>IN_0</name></connection>
<intersection>-4015 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-812,-4015,-770,-4015</points>
<connection>
<GID>1962</GID>
<name>OUT</name></connection>
<intersection>-812 0</intersection></hsegment></shape></wire>
<wire>
<ID>2224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795,-3903,-795,-3898</points>
<connection>
<GID>1911</GID>
<name>OUT_0</name></connection>
<intersection>-3903 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-796,-3908.5,-796,-3903</points>
<connection>
<GID>1922</GID>
<name>IN_1</name></connection>
<intersection>-3903 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-796,-3903,-795,-3903</points>
<intersection>-796 1</intersection>
<intersection>-795 0</intersection></hsegment></shape></wire>
<wire>
<ID>2225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-782,-3903,-782,-3897.5</points>
<connection>
<GID>1912</GID>
<name>OUT_0</name></connection>
<intersection>-3903 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-794,-3908.5,-794,-3903</points>
<connection>
<GID>1922</GID>
<name>IN_0</name></connection>
<intersection>-3903 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-794,-3903,-782,-3903</points>
<intersection>-794 1</intersection>
<intersection>-782 0</intersection></hsegment></shape></wire>
<wire>
<ID>2226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-831.5,-3923,-831.5,-3915.5</points>
<connection>
<GID>1914</GID>
<name>OUT</name></connection>
<intersection>-3923 9</intersection>
<intersection>-3918.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-818.5,-3931.5,-818.5,-3918.5</points>
<connection>
<GID>1924</GID>
<name>IN_1</name></connection>
<intersection>-3926.5 7</intersection>
<intersection>-3918.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-831.5,-3918.5,-818.5,-3918.5</points>
<intersection>-831.5 0</intersection>
<intersection>-818.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-818.5,-3926.5,-807,-3926.5</points>
<connection>
<GID>1943</GID>
<name>IN_0</name></connection>
<intersection>-818.5 1</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-885.5,-3923,-831.5,-3923</points>
<connection>
<GID>2065</GID>
<name>IN_0</name></connection>
<intersection>-831.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795,-3918,-795,-3914.5</points>
<connection>
<GID>1922</GID>
<name>OUT</name></connection>
<intersection>-3918 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-816.5,-3931.5,-816.5,-3918</points>
<connection>
<GID>1924</GID>
<name>IN_0</name></connection>
<intersection>-3928.5 6</intersection>
<intersection>-3925 8</intersection>
<intersection>-3918 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-816.5,-3918,-795,-3918</points>
<intersection>-816.5 1</intersection>
<intersection>-795 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-816.5,-3928.5,-807,-3928.5</points>
<connection>
<GID>1943</GID>
<name>IN_1</name></connection>
<intersection>-816.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-926,-3925,-816.5,-3925</points>
<connection>
<GID>2060</GID>
<name>IN_0</name></connection>
<intersection>-816.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-799.5,-4059,-799.5,-4006</points>
<connection>
<GID>2012</GID>
<name>IN_0</name></connection>
<intersection>-4006 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-799.5,-4006,-769.5,-4006</points>
<connection>
<GID>1964</GID>
<name>OUT</name></connection>
<intersection>-799.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-787,-4059,-787,-3998</points>
<connection>
<GID>2014</GID>
<name>IN_0</name></connection>
<intersection>-3998 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-787,-3998,-769,-3998</points>
<connection>
<GID>1966</GID>
<name>OUT</name></connection>
<intersection>-787 0</intersection></hsegment></shape></wire>
<wire>
<ID>2230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776,-4110.5,-776,-4110</points>
<intersection>-4110.5 1</intersection>
<intersection>-4110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-780,-4110.5,-776,-4110.5</points>
<connection>
<GID>1874</GID>
<name>OUT</name></connection>
<intersection>-776 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-776,-4110,-771.5,-4110</points>
<connection>
<GID>1968</GID>
<name>IN_0</name></connection>
<intersection>-776 0</intersection></hsegment></shape></wire>
<wire>
<ID>2231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-943.5,-3840.5,-884.5,-3840.5</points>
<connection>
<GID>1950</GID>
<name>OUT</name></connection>
<connection>
<GID>1940</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-861.5,-3876.5,-861.5,-3840.5</points>
<connection>
<GID>1930</GID>
<name>IN_1</name></connection>
<intersection>-3840.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-878.5,-3840.5,-861.5,-3840.5</points>
<connection>
<GID>1940</GID>
<name>Q</name></connection>
<intersection>-861.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-944,-3830.5,-897.5,-3830.5</points>
<connection>
<GID>1951</GID>
<name>OUT</name></connection>
<connection>
<GID>1941</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-848,-3876.5,-848,-3830.5</points>
<connection>
<GID>1931</GID>
<name>IN_1</name></connection>
<intersection>-3830.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-891.5,-3830.5,-848,-3830.5</points>
<connection>
<GID>1941</GID>
<name>Q</name></connection>
<intersection>-848 0</intersection></hsegment></shape></wire>
<wire>
<ID>2235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-945.5,-3819.5,-910.5,-3819.5</points>
<connection>
<GID>1952</GID>
<name>OUT</name></connection>
<connection>
<GID>1942</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-835,-3876.5,-835,-3819.5</points>
<connection>
<GID>1932</GID>
<name>IN_1</name></connection>
<intersection>-3819.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-904.5,-3819.5,-835,-3819.5</points>
<connection>
<GID>1942</GID>
<name>Q</name></connection>
<intersection>-835 0</intersection></hsegment></shape></wire>
<wire>
<ID>2237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-946,-3810.5,-918,-3810.5</points>
<connection>
<GID>1953</GID>
<name>OUT</name></connection>
<connection>
<GID>1944</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-822,-3876.5,-822,-3810.5</points>
<connection>
<GID>1933</GID>
<name>IN_1</name></connection>
<intersection>-3810.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-912,-3810.5,-822,-3810.5</points>
<connection>
<GID>1944</GID>
<name>Q</name></connection>
<intersection>-822 0</intersection></hsegment></shape></wire>
<wire>
<ID>2239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-947,-3803,-926.5,-3803</points>
<connection>
<GID>1954</GID>
<name>OUT</name></connection>
<connection>
<GID>1945</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-809.5,-3877,-809.5,-3803</points>
<connection>
<GID>1934</GID>
<name>IN_1</name></connection>
<intersection>-3803 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-920.5,-3803,-809.5,-3803</points>
<connection>
<GID>1945</GID>
<name>Q</name></connection>
<intersection>-809.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-948,-3795.5,-935.5,-3795.5</points>
<connection>
<GID>1955</GID>
<name>OUT</name></connection>
<connection>
<GID>1947</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-797,-3877,-797,-3795.5</points>
<connection>
<GID>1936</GID>
<name>IN_1</name></connection>
<intersection>-3795.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-929.5,-3795.5,-797,-3795.5</points>
<connection>
<GID>1947</GID>
<name>Q</name></connection>
<intersection>-797 0</intersection></hsegment></shape></wire>
<wire>
<ID>2243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-940.5,-3842.5,-940.5,-3791.5</points>
<connection>
<GID>1948</GID>
<name>OUT_0</name></connection>
<intersection>-3842.5 7</intersection>
<intersection>-3832.5 5</intersection>
<intersection>-3821.5 8</intersection>
<intersection>-3812.5 3</intersection>
<intersection>-3805 9</intersection>
<intersection>-3797.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-940.5,-3797.5,-935.5,-3797.5</points>
<connection>
<GID>1947</GID>
<name>clock</name></connection>
<intersection>-940.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-940.5,-3812.5,-918,-3812.5</points>
<connection>
<GID>1944</GID>
<name>clock</name></connection>
<intersection>-940.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-940.5,-3832.5,-897.5,-3832.5</points>
<connection>
<GID>1941</GID>
<name>clock</name></connection>
<intersection>-940.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-940.5,-3842.5,-884.5,-3842.5</points>
<connection>
<GID>1940</GID>
<name>clock</name></connection>
<intersection>-940.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-940.5,-3821.5,-910.5,-3821.5</points>
<connection>
<GID>1942</GID>
<name>clock</name></connection>
<intersection>-940.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-940.5,-3805,-926.5,-3805</points>
<connection>
<GID>1945</GID>
<name>clock</name></connection>
<intersection>-940.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-809.5,-4126.5,-809.5,-4119.5</points>
<connection>
<GID>2007</GID>
<name>OUT</name></connection>
<intersection>-4126.5 7</intersection>
<intersection>-4120 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-809.5,-4120,-608.5,-4120</points>
<intersection>-809.5 0</intersection>
<intersection>-771.5 5</intersection>
<intersection>-608.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-608.5,-4120,-608.5,-3636</points>
<connection>
<GID>1972</GID>
<name>IN_1</name></connection>
<intersection>-4120 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-771.5,-4120,-771.5,-4112</points>
<connection>
<GID>1968</GID>
<name>IN_1</name></connection>
<intersection>-4120 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-809.5,-4126.5,-797.5,-4126.5</points>
<connection>
<GID>1965</GID>
<name>J</name></connection>
<intersection>-809.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-765.5,-4106,-610.5,-4106</points>
<intersection>-765.5 11</intersection>
<intersection>-749 12</intersection>
<intersection>-610.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-610.5,-4106,-610.5,-3636</points>
<connection>
<GID>1972</GID>
<name>IN_0</name></connection>
<intersection>-4106 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-765.5,-4111,-765.5,-4106</points>
<connection>
<GID>1968</GID>
<name>OUT</name></connection>
<intersection>-4106 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-749,-4111,-749,-4106</points>
<connection>
<GID>1970</GID>
<name>N_in0</name></connection>
<intersection>-4106 1</intersection></vsegment></shape></wire>
<wire>
<ID>2246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-848.5,-4079.5,-848.5,-4074</points>
<connection>
<GID>2069</GID>
<name>clear</name></connection>
<intersection>-4079.5 1</intersection>
<intersection>-4074.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-916.5,-4079.5,-848.5,-4079.5</points>
<connection>
<GID>1871</GID>
<name>Q</name></connection>
<intersection>-848.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-848.5,-4074.5,-780.5,-4074.5</points>
<connection>
<GID>1997</GID>
<name>clear</name></connection>
<connection>
<GID>1996</GID>
<name>clear</name></connection>
<connection>
<GID>1995</GID>
<name>clear</name></connection>
<connection>
<GID>1994</GID>
<name>clear</name></connection>
<connection>
<GID>1993</GID>
<name>clear</name></connection>
<intersection>-848.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-919.5,-4300,-919.5,-4298</points>
<connection>
<GID>1897</GID>
<name>IN_0</name></connection>
<intersection>-4300 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-919.5,-4300,-915,-4300</points>
<connection>
<GID>1895</GID>
<name>OUT</name></connection>
<intersection>-919.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-919.5,-4294,-901.5,-4294</points>
<connection>
<GID>1897</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1892</GID>
<name>clear</name></connection>
<intersection>-919.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-919.5,-4294,-919.5,-4288</points>
<intersection>-4294 1</intersection>
<intersection>-4288 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-919.5,-4288,-904.5,-4288</points>
<connection>
<GID>1892</GID>
<name>J</name></connection>
<intersection>-919.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2249</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-898.5,-4292,-895.5,-4292</points>
<connection>
<GID>1892</GID>
<name>nQ</name></connection>
<connection>
<GID>1898</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-909,-4299,-874.5,-4299</points>
<connection>
<GID>1895</GID>
<name>IN_1</name></connection>
<intersection>-874.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-874.5,-4299,-874.5,-4298</points>
<connection>
<GID>1901</GID>
<name>OUT</name></connection>
<intersection>-4299 1</intersection></vsegment></shape></wire>
<wire>
<ID>2251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-838,-4288,-838,-4273</points>
<connection>
<GID>2153</GID>
<name>clear</name></connection>
<intersection>-4288 1</intersection>
<intersection>-4273.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-898.5,-4288,-838,-4288</points>
<connection>
<GID>1892</GID>
<name>Q</name></connection>
<intersection>-838 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-838,-4273.5,-770,-4273.5</points>
<connection>
<GID>2076</GID>
<name>clear</name></connection>
<connection>
<GID>2075</GID>
<name>clear</name></connection>
<connection>
<GID>2073</GID>
<name>clear</name></connection>
<connection>
<GID>2072</GID>
<name>clear</name></connection>
<connection>
<GID>2070</GID>
<name>clear</name></connection>
<intersection>-838 0</intersection></hsegment></shape></wire>
<wire>
<ID>2252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-921,-4523,-921,-4521</points>
<connection>
<GID>1937</GID>
<name>IN_0</name></connection>
<intersection>-4523 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-921,-4523,-916.5,-4523</points>
<connection>
<GID>1906</GID>
<name>OUT</name></connection>
<intersection>-921 0</intersection></hsegment></shape></wire>
<wire>
<ID>2253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-921,-4517,-903,-4517</points>
<connection>
<GID>1937</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1903</GID>
<name>clear</name></connection>
<intersection>-921 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-921,-4517,-921,-4511</points>
<intersection>-4517 1</intersection>
<intersection>-4511 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-921,-4511,-906,-4511</points>
<connection>
<GID>1903</GID>
<name>J</name></connection>
<intersection>-921 3</intersection></hsegment></shape></wire>
<wire>
<ID>2254</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-900,-4515,-897,-4515</points>
<connection>
<GID>1903</GID>
<name>nQ</name></connection>
<connection>
<GID>1957</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-910.5,-4522,-876,-4522</points>
<connection>
<GID>1906</GID>
<name>IN_1</name></connection>
<intersection>-876 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-876,-4522,-876,-4521</points>
<connection>
<GID>1960</GID>
<name>OUT</name></connection>
<intersection>-4522 1</intersection></vsegment></shape></wire>
<wire>
<ID>2256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-844.5,-4511,-844.5,-4495</points>
<connection>
<GID>2401</GID>
<name>clear</name></connection>
<intersection>-4511 1</intersection>
<intersection>-4495.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-900,-4511,-844.5,-4511</points>
<connection>
<GID>1903</GID>
<name>Q</name></connection>
<intersection>-844.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-844.5,-4495.5,-776.5,-4495.5</points>
<connection>
<GID>2169</GID>
<name>clear</name></connection>
<connection>
<GID>2158</GID>
<name>clear</name></connection>
<connection>
<GID>2157</GID>
<name>clear</name></connection>
<connection>
<GID>2156</GID>
<name>clear</name></connection>
<connection>
<GID>2155</GID>
<name>clear</name></connection>
<intersection>-844.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-919,-4756.5,-919,-4754.5</points>
<connection>
<GID>1971</GID>
<name>IN_0</name></connection>
<intersection>-4756.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-919,-4756.5,-914.5,-4756.5</points>
<connection>
<GID>1967</GID>
<name>OUT</name></connection>
<intersection>-919 0</intersection></hsegment></shape></wire>
<wire>
<ID>2258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-919,-4750.5,-901,-4750.5</points>
<connection>
<GID>1971</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1963</GID>
<name>clear</name></connection>
<intersection>-919 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-919,-4750.5,-919,-4744.5</points>
<intersection>-4750.5 1</intersection>
<intersection>-4744.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-919,-4744.5,-904,-4744.5</points>
<connection>
<GID>1963</GID>
<name>J</name></connection>
<intersection>-919 3</intersection></hsegment></shape></wire>
<wire>
<ID>2259</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-898,-4748.5,-895,-4748.5</points>
<connection>
<GID>1963</GID>
<name>nQ</name></connection>
<connection>
<GID>1974</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-908.5,-4755.5,-874,-4755.5</points>
<connection>
<GID>1967</GID>
<name>IN_1</name></connection>
<intersection>-874 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-874,-4755.5,-874,-4754.5</points>
<connection>
<GID>1977</GID>
<name>OUT</name></connection>
<intersection>-4755.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-842.5,-4744.5,-842.5,-4729</points>
<connection>
<GID>2440</GID>
<name>clear</name></connection>
<intersection>-4744.5 1</intersection>
<intersection>-4729.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-898,-4744.5,-842.5,-4744.5</points>
<connection>
<GID>1963</GID>
<name>Q</name></connection>
<intersection>-842.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-842.5,-4729.5,-774.5,-4729.5</points>
<connection>
<GID>2406</GID>
<name>clear</name></connection>
<connection>
<GID>2405</GID>
<name>clear</name></connection>
<connection>
<GID>2404</GID>
<name>clear</name></connection>
<connection>
<GID>2403</GID>
<name>clear</name></connection>
<connection>
<GID>2402</GID>
<name>clear</name></connection>
<intersection>-842.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-896.5,-4985,-896.5,-4983</points>
<connection>
<GID>1983</GID>
<name>IN_0</name></connection>
<intersection>-4985 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-896.5,-4985,-892,-4985</points>
<connection>
<GID>1981</GID>
<name>OUT</name></connection>
<intersection>-896.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-896.5,-4979,-878.5,-4979</points>
<connection>
<GID>1983</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1979</GID>
<name>clear</name></connection>
<intersection>-896.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-896.5,-4979,-896.5,-4973</points>
<intersection>-4979 1</intersection>
<intersection>-4973 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-896.5,-4973,-881.5,-4973</points>
<connection>
<GID>1979</GID>
<name>J</name></connection>
<intersection>-896.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2264</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-875.5,-4977,-872.5,-4977</points>
<connection>
<GID>1979</GID>
<name>nQ</name></connection>
<connection>
<GID>1985</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-790,-4137,-790,-4126.5</points>
<intersection>-4137 2</intersection>
<intersection>-4126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-791.5,-4126.5,-790,-4126.5</points>
<connection>
<GID>1965</GID>
<name>Q</name></connection>
<intersection>-790 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-790,-4137,-788,-4137</points>
<connection>
<GID>1969</GID>
<name>IN_0</name></connection>
<intersection>-790 0</intersection></hsegment></shape></wire>
<wire>
<ID>2266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-841,-4257.5,-841,-4209.5</points>
<connection>
<GID>2107</GID>
<name>IN_0</name></connection>
<intersection>-4209.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-841,-4209.5,-768.5,-4209.5</points>
<connection>
<GID>1973</GID>
<name>OUT</name></connection>
<intersection>-841 0</intersection></hsegment></shape></wire>
<wire>
<ID>2267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-760.5,-4208.5,-760.5,-4138</points>
<intersection>-4208.5 2</intersection>
<intersection>-4161.5 3</intersection>
<intersection>-4138 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-782,-4138,-760.5,-4138</points>
<connection>
<GID>1969</GID>
<name>OUT</name></connection>
<intersection>-760.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-762.5,-4208.5,-760.5,-4208.5</points>
<connection>
<GID>1973</GID>
<name>IN_1</name></connection>
<intersection>-760.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-760.5,-4161.5,-743,-4161.5</points>
<intersection>-760.5 0</intersection>
<intersection>-748 9</intersection>
<intersection>-743 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-743,-4200,-743,-4161.5</points>
<intersection>-4200 5</intersection>
<intersection>-4190 6</intersection>
<intersection>-4183 7</intersection>
<intersection>-4173.5 8</intersection>
<intersection>-4161.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-750.5,-4200,-743,-4200</points>
<connection>
<GID>1975</GID>
<name>IN_1</name></connection>
<intersection>-743 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-750.5,-4190,-743,-4190</points>
<connection>
<GID>1976</GID>
<name>IN_1</name></connection>
<intersection>-743 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-749,-4183,-743,-4183</points>
<connection>
<GID>1978</GID>
<name>IN_1</name></connection>
<intersection>-743 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-748.5,-4173.5,-743,-4173.5</points>
<connection>
<GID>1980</GID>
<name>IN_1</name></connection>
<intersection>-743 4</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-748,-4166.5,-748,-4161.5</points>
<connection>
<GID>1982</GID>
<name>IN_1</name></connection>
<intersection>-4161.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>2268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-827.5,-4257.5,-827.5,-4198</points>
<connection>
<GID>2110</GID>
<name>IN_0</name></connection>
<intersection>-4198 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-827.5,-4198,-756.5,-4198</points>
<intersection>-827.5 0</intersection>
<intersection>-756.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-756.5,-4201,-756.5,-4198</points>
<connection>
<GID>1975</GID>
<name>OUT</name></connection>
<intersection>-4198 1</intersection></vsegment></shape></wire>
<wire>
<ID>2269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-814.5,-4257.5,-814.5,-4189.5</points>
<connection>
<GID>2112</GID>
<name>IN_0</name></connection>
<intersection>-4189.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-814.5,-4189.5,-756.5,-4189.5</points>
<intersection>-814.5 0</intersection>
<intersection>-756.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-756.5,-4191,-756.5,-4189.5</points>
<connection>
<GID>1976</GID>
<name>OUT</name></connection>
<intersection>-4189.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-801.5,-4257.5,-801.5,-4182</points>
<connection>
<GID>2114</GID>
<name>IN_0</name></connection>
<intersection>-4182 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-801.5,-4182,-755,-4182</points>
<intersection>-801.5 0</intersection>
<intersection>-755 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-755,-4184,-755,-4182</points>
<connection>
<GID>1978</GID>
<name>OUT</name></connection>
<intersection>-4182 1</intersection></vsegment></shape></wire>
<wire>
<ID>2271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-789,-4258,-789,-4174.5</points>
<connection>
<GID>2116</GID>
<name>IN_0</name></connection>
<intersection>-4174.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-789,-4174.5,-754.5,-4174.5</points>
<connection>
<GID>1980</GID>
<name>OUT</name></connection>
<intersection>-789 0</intersection></hsegment></shape></wire>
<wire>
<ID>2272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-776.5,-4258,-776.5,-4167.5</points>
<connection>
<GID>2120</GID>
<name>IN_0</name></connection>
<intersection>-4167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-776.5,-4167.5,-754,-4167.5</points>
<connection>
<GID>1982</GID>
<name>OUT</name></connection>
<intersection>-776.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-769.5,-4309.5,-769.5,-4309</points>
<intersection>-4309.5 1</intersection>
<intersection>-4309 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-772,-4309.5,-769.5,-4309.5</points>
<connection>
<GID>1876</GID>
<name>OUT</name></connection>
<intersection>-769.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-769.5,-4309,-766.5,-4309</points>
<connection>
<GID>1984</GID>
<name>IN_0</name></connection>
<intersection>-769.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-799,-4323,-799,-4318.5</points>
<connection>
<GID>2103</GID>
<name>OUT</name></connection>
<intersection>-4323 7</intersection>
<intersection>-4319 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-799,-4319,-593.5,-4319</points>
<intersection>-799 0</intersection>
<intersection>-766.5 5</intersection>
<intersection>-593.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-593.5,-4319,-593.5,-3636.5</points>
<connection>
<GID>1987</GID>
<name>IN_1</name></connection>
<intersection>-4319 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-766.5,-4319,-766.5,-4311</points>
<connection>
<GID>1984</GID>
<name>IN_1</name></connection>
<intersection>-4319 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-799,-4323,-789.5,-4323</points>
<connection>
<GID>1989</GID>
<name>J</name></connection>
<intersection>-799 0</intersection></hsegment></shape></wire>
<wire>
<ID>2275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-755.5,-4310,-755.5,-4309.5</points>
<intersection>-4310 2</intersection>
<intersection>-4309.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-755.5,-4309.5,-595.5,-4309.5</points>
<connection>
<GID>1986</GID>
<name>N_in0</name></connection>
<intersection>-755.5 0</intersection>
<intersection>-595.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-760.5,-4310,-755.5,-4310</points>
<connection>
<GID>1984</GID>
<name>OUT</name></connection>
<intersection>-755.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-595.5,-4309.5,-595.5,-3636.5</points>
<connection>
<GID>1987</GID>
<name>IN_0</name></connection>
<intersection>-4309.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-779.5,-4332.5,-779.5,-4323</points>
<intersection>-4332.5 2</intersection>
<intersection>-4323 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-783.5,-4323,-779.5,-4323</points>
<connection>
<GID>1989</GID>
<name>Q</name></connection>
<intersection>-779.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-779.5,-4332.5,-775,-4332.5</points>
<connection>
<GID>1990</GID>
<name>IN_0</name></connection>
<intersection>-779.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-770.5,-4467,-770.5,-4333.5</points>
<intersection>-4467 2</intersection>
<intersection>-4409.5 3</intersection>
<intersection>-4333.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-770.5,-4333.5,-769,-4333.5</points>
<connection>
<GID>1990</GID>
<name>OUT</name></connection>
<intersection>-770.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-771.5,-4467,-770.5,-4467</points>
<connection>
<GID>1991</GID>
<name>IN_1</name></connection>
<intersection>-770.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-770.5,-4409.5,-751.5,-4409.5</points>
<intersection>-770.5 0</intersection>
<intersection>-751.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-751.5,-4461,-751.5,-4409.5</points>
<intersection>-4461 5</intersection>
<intersection>-4451.5 6</intersection>
<intersection>-4442 7</intersection>
<intersection>-4433.5 8</intersection>
<intersection>-4425 9</intersection>
<intersection>-4409.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-760.5,-4461,-751.5,-4461</points>
<connection>
<GID>1992</GID>
<name>IN_1</name></connection>
<intersection>-751.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-760.5,-4451.5,-751.5,-4451.5</points>
<connection>
<GID>2013</GID>
<name>IN_1</name></connection>
<intersection>-751.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-759.5,-4442,-751.5,-4442</points>
<connection>
<GID>2016</GID>
<name>IN_1</name></connection>
<intersection>-751.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-759,-4433.5,-751.5,-4433.5</points>
<connection>
<GID>2029</GID>
<name>IN_1</name></connection>
<intersection>-751.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-758,-4425,-751.5,-4425</points>
<connection>
<GID>2030</GID>
<name>IN_1</name></connection>
<intersection>-751.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-847.5,-4479.5,-847.5,-4468</points>
<connection>
<GID>2352</GID>
<name>IN_0</name></connection>
<intersection>-4468 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-847.5,-4468,-777.5,-4468</points>
<connection>
<GID>1991</GID>
<name>OUT</name></connection>
<intersection>-847.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-972.5,-4111.5,-972.5,-3948</points>
<intersection>-4111.5 13</intersection>
<intersection>-4021.5 1</intersection>
<intersection>-4011.5 3</intersection>
<intersection>-4000.5 5</intersection>
<intersection>-3991.5 7</intersection>
<intersection>-3984 9</intersection>
<intersection>-3976.5 11</intersection>
<intersection>-3955.5 16</intersection>
<intersection>-3948 15</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-972.5,-4021.5,-941.5,-4021.5</points>
<connection>
<GID>2025</GID>
<name>IN_0</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-972.5,-4011.5,-942,-4011.5</points>
<connection>
<GID>2026</GID>
<name>IN_0</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-972.5,-4000.5,-943.5,-4000.5</points>
<connection>
<GID>2027</GID>
<name>IN_0</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-972.5,-3991.5,-944,-3991.5</points>
<connection>
<GID>2028</GID>
<name>IN_0</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-972.5,-3984,-945,-3984</points>
<connection>
<GID>2039</GID>
<name>IN_0</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-972.5,-3976.5,-946,-3976.5</points>
<connection>
<GID>2067</GID>
<name>IN_0</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-972.5,-4111.5,-786,-4111.5</points>
<connection>
<GID>1874</GID>
<name>IN_1</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-972.5,-3948,-786,-3948</points>
<connection>
<GID>1935</GID>
<name>IN_1</name></connection>
<intersection>-972.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-980.5,-3955.5,-972.5,-3955.5</points>
<intersection>-980.5 17</intersection>
<intersection>-972.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-980.5,-3955.5,-980.5,-3955</points>
<connection>
<GID>2089</GID>
<name>OUT</name></connection>
<intersection>-3955.5 16</intersection></vsegment></shape></wire>
<wire>
<ID>2280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-852.5,-4068,-852.5,-4064.5</points>
<connection>
<GID>2008</GID>
<name>OUT</name></connection>
<intersection>-4068 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-852.5,-4068,-851.5,-4068</points>
<connection>
<GID>2069</GID>
<name>IN_0</name></connection>
<intersection>-852.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-839,-4068.5,-839,-4064.5</points>
<connection>
<GID>2009</GID>
<name>OUT</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-839,-4068.5,-835.5,-4068.5</points>
<connection>
<GID>1993</GID>
<name>IN_0</name></connection>
<intersection>-839 0</intersection></hsegment></shape></wire>
<wire>
<ID>2282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-826,-4068.5,-826,-4064.5</points>
<connection>
<GID>2010</GID>
<name>OUT</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-826,-4068.5,-822,-4068.5</points>
<connection>
<GID>1994</GID>
<name>IN_0</name></connection>
<intersection>-826 0</intersection></hsegment></shape></wire>
<wire>
<ID>2283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-810,-4068.5,-810,-4064.5</points>
<intersection>-4068.5 1</intersection>
<intersection>-4064.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-810,-4068.5,-807,-4068.5</points>
<connection>
<GID>1995</GID>
<name>IN_0</name></connection>
<intersection>-810 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-813,-4064.5,-810,-4064.5</points>
<connection>
<GID>2011</GID>
<name>OUT</name></connection>
<intersection>-810 0</intersection></hsegment></shape></wire>
<wire>
<ID>2284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-800.5,-4067,-800.5,-4065</points>
<connection>
<GID>2012</GID>
<name>OUT</name></connection>
<intersection>-4067 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-800.5,-4067,-796.5,-4067</points>
<intersection>-800.5 0</intersection>
<intersection>-796.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-796.5,-4068.5,-796.5,-4067</points>
<connection>
<GID>1996</GID>
<name>IN_0</name></connection>
<intersection>-4067 1</intersection></vsegment></shape></wire>
<wire>
<ID>2285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-788,-4067,-788,-4065</points>
<connection>
<GID>2014</GID>
<name>OUT</name></connection>
<intersection>-4067 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-788,-4067,-783.5,-4067</points>
<intersection>-788 0</intersection>
<intersection>-783.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-783.5,-4068.5,-783.5,-4067</points>
<connection>
<GID>1997</GID>
<name>IN_0</name></connection>
<intersection>-4067 1</intersection></vsegment></shape></wire>
<wire>
<ID>2286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-841.5,-4076,-841.5,-4068</points>
<connection>
<GID>1998</GID>
<name>IN_0</name></connection>
<intersection>-4068 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-845.5,-4068,-841.5,-4068</points>
<connection>
<GID>2069</GID>
<name>OUT_0</name></connection>
<intersection>-841.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-826.5,-4076,-826.5,-4068.5</points>
<connection>
<GID>1999</GID>
<name>IN_0</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-829.5,-4068.5,-826.5,-4068.5</points>
<connection>
<GID>1993</GID>
<name>OUT_0</name></connection>
<intersection>-826.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-811.5,-4076,-811.5,-4068.5</points>
<connection>
<GID>2000</GID>
<name>IN_0</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-816,-4068.5,-811.5,-4068.5</points>
<connection>
<GID>1994</GID>
<name>OUT_0</name></connection>
<intersection>-811.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-800,-4075.5,-800,-4068.5</points>
<connection>
<GID>2001</GID>
<name>IN_0</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-801,-4068.5,-800,-4068.5</points>
<connection>
<GID>1995</GID>
<name>OUT_0</name></connection>
<intersection>-800 0</intersection></hsegment></shape></wire>
<wire>
<ID>2290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-787,-4076,-787,-4068.5</points>
<connection>
<GID>2002</GID>
<name>IN_0</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-790.5,-4068.5,-787,-4068.5</points>
<connection>
<GID>1996</GID>
<name>OUT_0</name></connection>
<intersection>-787 0</intersection></hsegment></shape></wire>
<wire>
<ID>2291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-774,-4075.5,-774,-4068.5</points>
<connection>
<GID>2003</GID>
<name>IN_0</name></connection>
<intersection>-4068.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-777.5,-4068.5,-774,-4068.5</points>
<connection>
<GID>1997</GID>
<name>OUT_0</name></connection>
<intersection>-774 0</intersection></hsegment></shape></wire>
<wire>
<ID>2292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-841.5,-4085.5,-841.5,-4080</points>
<connection>
<GID>1998</GID>
<name>OUT_0</name></connection>
<intersection>-4085.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-826.5,-4091.5,-826.5,-4085.5</points>
<connection>
<GID>2004</GID>
<name>IN_3</name></connection>
<intersection>-4085.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-841.5,-4085.5,-826.5,-4085.5</points>
<intersection>-841.5 0</intersection>
<intersection>-826.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-826.5,-4085,-826.5,-4080</points>
<connection>
<GID>1999</GID>
<name>OUT_0</name></connection>
<intersection>-4085 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-824.5,-4091.5,-824.5,-4085</points>
<connection>
<GID>2004</GID>
<name>IN_2</name></connection>
<intersection>-4085 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-826.5,-4085,-824.5,-4085</points>
<intersection>-826.5 0</intersection>
<intersection>-824.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-811.5,-4085.5,-811.5,-4080</points>
<connection>
<GID>2000</GID>
<name>OUT_0</name></connection>
<intersection>-4085.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-822.5,-4091.5,-822.5,-4085.5</points>
<connection>
<GID>2004</GID>
<name>IN_1</name></connection>
<intersection>-4085.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-822.5,-4085.5,-811.5,-4085.5</points>
<intersection>-822.5 1</intersection>
<intersection>-811.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-800,-4086.5,-800,-4079.5</points>
<connection>
<GID>2001</GID>
<name>OUT_0</name></connection>
<intersection>-4086.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-820.5,-4091.5,-820.5,-4086.5</points>
<connection>
<GID>2004</GID>
<name>IN_0</name></connection>
<intersection>-4086.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-820.5,-4086.5,-800,-4086.5</points>
<intersection>-820.5 1</intersection>
<intersection>-800 0</intersection></hsegment></shape></wire>
<wire>
<ID>2296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-787,-4085,-787,-4080</points>
<connection>
<GID>2002</GID>
<name>OUT_0</name></connection>
<intersection>-4085 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-788,-4090.5,-788,-4085</points>
<connection>
<GID>2006</GID>
<name>IN_1</name></connection>
<intersection>-4085 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-788,-4085,-787,-4085</points>
<intersection>-788 1</intersection>
<intersection>-787 0</intersection></hsegment></shape></wire>
<wire>
<ID>2297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-774,-4085,-774,-4079.5</points>
<connection>
<GID>2003</GID>
<name>OUT_0</name></connection>
<intersection>-4085 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-786,-4090.5,-786,-4085</points>
<connection>
<GID>2006</GID>
<name>IN_0</name></connection>
<intersection>-4085 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-786,-4085,-774,-4085</points>
<intersection>-786 1</intersection>
<intersection>-774 0</intersection></hsegment></shape></wire>
<wire>
<ID>2298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-823.5,-4100.5,-823.5,-4097.5</points>
<connection>
<GID>2004</GID>
<name>OUT</name></connection>
<intersection>-4100.5 2</intersection>
<intersection>-4098 8</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-810.5,-4113.5,-810.5,-4100.5</points>
<connection>
<GID>2007</GID>
<name>IN_1</name></connection>
<intersection>-4108.5 7</intersection>
<intersection>-4100.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-823.5,-4100.5,-810.5,-4100.5</points>
<intersection>-823.5 0</intersection>
<intersection>-810.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-810.5,-4108.5,-799,-4108.5</points>
<connection>
<GID>2020</GID>
<name>IN_0</name></connection>
<intersection>-810.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-886.5,-4098,-823.5,-4098</points>
<intersection>-886.5 9</intersection>
<intersection>-823.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-886.5,-4098,-886.5,-4090.5</points>
<connection>
<GID>1888</GID>
<name>IN_0</name></connection>
<intersection>-4098 8</intersection></vsegment></shape></wire>
<wire>
<ID>2299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-834,-4479.5,-834,-4462</points>
<connection>
<GID>2354</GID>
<name>IN_0</name></connection>
<intersection>-4462 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-834,-4462,-766.5,-4462</points>
<connection>
<GID>1992</GID>
<name>OUT</name></connection>
<intersection>-834 0</intersection></hsegment></shape></wire>
<wire>
<ID>2300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-821,-4479.5,-821,-4452.5</points>
<connection>
<GID>2356</GID>
<name>IN_0</name></connection>
<intersection>-4452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-821,-4452.5,-766.5,-4452.5</points>
<connection>
<GID>2013</GID>
<name>OUT</name></connection>
<intersection>-821 0</intersection></hsegment></shape></wire>
<wire>
<ID>2301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808,-4479.5,-808,-4443</points>
<connection>
<GID>2357</GID>
<name>IN_0</name></connection>
<intersection>-4443 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-808,-4443,-765.5,-4443</points>
<connection>
<GID>2016</GID>
<name>OUT</name></connection>
<intersection>-808 0</intersection></hsegment></shape></wire>
<wire>
<ID>2302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-795.5,-4480,-795.5,-4434.5</points>
<connection>
<GID>2358</GID>
<name>IN_0</name></connection>
<intersection>-4434.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-795.5,-4434.5,-765,-4434.5</points>
<connection>
<GID>2029</GID>
<name>OUT</name></connection>
<intersection>-795.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-787,-4100,-787,-4096.5</points>
<connection>
<GID>2006</GID>
<name>OUT</name></connection>
<intersection>-4100 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-808.5,-4113.5,-808.5,-4100</points>
<connection>
<GID>2007</GID>
<name>IN_0</name></connection>
<intersection>-4110.5 6</intersection>
<intersection>-4104 7</intersection>
<intersection>-4100 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-808.5,-4100,-787,-4100</points>
<intersection>-808.5 1</intersection>
<intersection>-787 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-808.5,-4110.5,-799,-4110.5</points>
<connection>
<GID>2020</GID>
<name>IN_1</name></connection>
<intersection>-808.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-927,-4104,-808.5,-4104</points>
<intersection>-927 8</intersection>
<intersection>-808.5 1</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-927,-4104,-927,-4092.5</points>
<connection>
<GID>1872</GID>
<name>IN_0</name></connection>
<intersection>-4104 7</intersection></vsegment></shape></wire>
<wire>
<ID>2304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-783,-4480,-783,-4426</points>
<connection>
<GID>2359</GID>
<name>IN_0</name></connection>
<intersection>-4426 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-783,-4426,-764,-4426</points>
<connection>
<GID>2030</GID>
<name>OUT</name></connection>
<intersection>-783 0</intersection></hsegment></shape></wire>
<wire>
<ID>2305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-776.5,-4531.5,-770,-4531.5</points>
<connection>
<GID>1880</GID>
<name>OUT</name></connection>
<connection>
<GID>2031</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-805.5,-4548,-805.5,-4540.5</points>
<connection>
<GID>2345</GID>
<name>OUT</name></connection>
<intersection>-4548 4</intersection>
<intersection>-4541.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-805.5,-4541.5,-579.5,-4541.5</points>
<intersection>-805.5 0</intersection>
<intersection>-770 7</intersection>
<intersection>-579.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-579.5,-4541.5,-579.5,-3636.5</points>
<connection>
<GID>2051</GID>
<name>IN_1</name></connection>
<intersection>-4541.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-805.5,-4548,-795,-4548</points>
<connection>
<GID>2033</GID>
<name>J</name></connection>
<intersection>-805.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-770,-4541.5,-770,-4533.5</points>
<connection>
<GID>2031</GID>
<name>IN_1</name></connection>
<intersection>-4541.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-162.075,90.9046,324.525,-149.613</PageViewport>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>19,31</position>
<gparam>LABEL_TEXT Default Power</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>-69.5,39.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>299 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>19</ID>
<type>BB_CLOCK</type>
<position>-84,32.5</position>
<output>
<ID>CLK</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>48,-97.5</position>
<gparam>LABEL_TEXT Checking condition for 60</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>-83.5,41.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>249.5,-16.5</position>
<gparam>LABEL_TEXT Problematic Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>BA_NAND4</type>
<position>226.5,38.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>61 </input>
<input>
<ID>IN_3</ID>67 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_DFF_LOW</type>
<position>27.5,-31.5</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>58</ID>
<type>BE_JKFF_LOW_NT</type>
<position>9.5,13</position>
<input>
<ID>J</ID>92 </input>
<input>
<ID>K</ID>98 </input>
<output>
<ID>Q</ID>34 </output>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>66 </input>
<output>
<ID>nQ</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>60</ID>
<type>BE_JKFF_LOW_NT</type>
<position>59,12.5</position>
<input>
<ID>J</ID>133 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>39 </output>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>66 </input>
<output>
<ID>nQ</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_DFF_LOW</type>
<position>70.5,-31</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>63</ID>
<type>BE_JKFF_LOW_NT</type>
<position>85,13</position>
<input>
<ID>J</ID>135 </input>
<input>
<ID>K</ID>136 </input>
<output>
<ID>Q</ID>45 </output>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>66 </input>
<output>
<ID>nQ</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>65</ID>
<type>BE_JKFF_LOW_NT</type>
<position>115,12.5</position>
<input>
<ID>J</ID>137 </input>
<input>
<ID>K</ID>138 </input>
<output>
<ID>Q</ID>50 </output>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>66 </input>
<output>
<ID>nQ</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>BE_JKFF_LOW_NT</type>
<position>153.5,10.5</position>
<input>
<ID>J</ID>139 </input>
<input>
<ID>K</ID>140 </input>
<output>
<ID>Q</ID>61 </output>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>66 </input>
<output>
<ID>nQ</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>BE_JKFF_LOW_NT</type>
<position>202,10</position>
<input>
<ID>J</ID>141 </input>
<input>
<ID>K</ID>142 </input>
<output>
<ID>Q</ID>67 </output>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_DFF_LOW</type>
<position>100,-31</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>26,22</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>25,4.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>419 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_AND2</type>
<position>67,22</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>69.5,3.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_AND2</type>
<position>96.5,20.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND2</type>
<position>99,2</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>123,19.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>124.5,2</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>170,20.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND2</type>
<position>170.5,3</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_DFF_LOW</type>
<position>128.5,-31</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>71 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_OR2</type>
<position>40,12.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_DFF_LOW</type>
<position>174.5,-31</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR2</type>
<position>76.5,13.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_OR2</type>
<position>105,13</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_OR2</type>
<position>134,12.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_OR2</type>
<position>178,12</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_DFF_LOW</type>
<position>222.5,-31.5</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>109</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>226.5,-11</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>45 </input>
<input>
<ID>IN_3</ID>50 </input>
<input>
<ID>IN_4</ID>61 </input>
<input>
<ID>IN_5</ID>67 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>496</ID>
<type>AE_DFF_LOW</type>
<position>-54,4.5</position>
<input>
<ID>IN_0</ID>417 </input>
<output>
<ID>OUTINV_0</ID>419 </output>
<output>
<ID>OUT_0</ID>418 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>497</ID>
<type>CC_PULSE</type>
<position>-100,9.5</position>
<output>
<ID>OUT_0</ID>414 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>246,-41.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<input>
<ID>IN_4</ID>73 </input>
<input>
<ID>IN_5</ID>74 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>498</ID>
<type>CC_PULSE</type>
<position>-100,-8</position>
<output>
<ID>OUT_0</ID>412 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>EE_VDD</type>
<position>-49.5,45</position>
<output>
<ID>OUT_0</ID>300 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>501</ID>
<type>AE_OR2</type>
<position>-63,-7</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>412 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>AE_SMALL_INVERTER</type>
<position>-80.5,9.5</position>
<input>
<ID>IN_0</ID>414 </input>
<output>
<ID>OUT_0</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>43.5,-82</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>AI_XOR2</type>
<position>-66,5.5</position>
<input>
<ID>IN_0</ID>412 </input>
<input>
<ID>IN_1</ID>415 </input>
<output>
<ID>OUT</ID>417 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_LABEL</type>
<position>-96,16</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>117.5,-68.5</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_LABEL</type>
<position>-97,-13</position>
<gparam>LABEL_TEXT Text</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_AND2</type>
<position>180.5,-67</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AI_XOR2</type>
<position>-6,24</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>AI_XOR2</type>
<position>45,26.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AI_XOR2</type>
<position>81.5,27</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AI_XOR2</type>
<position>110,26.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AI_XOR2</type>
<position>140,26.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AI_XOR2</type>
<position>187.5,28.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_AND4</type>
<position>22,-104</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>129 </input>
<input>
<ID>IN_2</ID>126 </input>
<input>
<ID>IN_3</ID>419 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_INVERTER</type>
<position>37.5,-59</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_INVERTER</type>
<position>50,-60</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_INVERTER</type>
<position>114,-59</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_INVERTER</type>
<position>121,-59</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_INVERTER</type>
<position>178.5,-58.5</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_INVERTER</type>
<position>184,-58</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>246,-51.5</position>
<gparam>LABEL_TEXT Actual Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>-32.5,-14.5</position>
<gparam>LABEL_TEXT Clock input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>360</ID>
<type>AA_AND2</type>
<position>-56.5,38.5</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>299 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>72.5,48</position>
<gparam>LABEL_TEXT Setting Mode</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_LABEL</type>
<position>-77.5,49</position>
<gparam>LABEL_TEXT On/Off- Settings/Cycle</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>AA_LABEL</type>
<position>-33,17</position>
<gparam>LABEL_TEXT Direction</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-81.5,41.5,-72.5,41.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76,32.5,-76,38.5</points>
<intersection>32.5 2</intersection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,38.5,-72.5,38.5</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>-76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80,32.5,-76,32.5</points>
<connection>
<GID>19</GID>
<name>CLK</name></connection>
<intersection>-76 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-17,234.5,38.5</points>
<intersection>-17 2</intersection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,38.5,234.5,38.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-17,234.5,-17</points>
<intersection>9.5 15</intersection>
<intersection>59 14</intersection>
<intersection>85 10</intersection>
<intersection>115 18</intersection>
<intersection>153.5 16</intersection>
<intersection>202 17</intersection>
<intersection>234.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>85,-17,85,9</points>
<connection>
<GID>63</GID>
<name>clear</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>59,-17,59,8.5</points>
<connection>
<GID>60</GID>
<name>clear</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>9.5,-17,9.5,9</points>
<connection>
<GID>58</GID>
<name>clear</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>153.5,-17,153.5,6.5</points>
<connection>
<GID>67</GID>
<name>clear</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>202,-17,202,6</points>
<connection>
<GID>69</GID>
<name>clear</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>115,-17,115,8.5</points>
<connection>
<GID>65</GID>
<name>clear</name></connection>
<intersection>-17 2</intersection></vsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,-8,-70.5,17</points>
<intersection>-8 1</intersection>
<intersection>17 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98,-8,-66,-8</points>
<connection>
<GID>501</GID>
<name>IN_1</name></connection>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-70.5,17,-65,17</points>
<intersection>-70.5 0</intersection>
<intersection>-65 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-65,8.5,-65,17</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>17 4</intersection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-6,-84,9.5</points>
<intersection>-6 3</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98,9.5,-82.5,9.5</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-84,-6,-66,-6</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>-84 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,8.5,-67,9.5</points>
<connection>
<GID>504</GID>
<name>IN_1</name></connection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78.5,9.5,-67,9.5</points>
<connection>
<GID>502</GID>
<name>OUT_0</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-66,2,-60.5,2</points>
<intersection>-66 5</intersection>
<intersection>-60.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-60.5,2,-60.5,6.5</points>
<intersection>2 1</intersection>
<intersection>6.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-66,2,-66,2.5</points>
<connection>
<GID>504</GID>
<name>OUT</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-60.5,6.5,-57,6.5</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>-60.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,6.5,-46.5,23</points>
<intersection>6.5 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51,6.5,-46.5,6.5</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46.5,23,23,23</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,3.5,22,3.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<connection>
<GID>496</GID>
<name>OUTINV_0</name></connection>
<intersection>-21.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-21.5,-101,-21.5,3.5</points>
<intersection>-101 8</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-21.5,-101,19,-101</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>-21.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-29.5,18.5,21</points>
<intersection>-29.5 8</intersection>
<intersection>-23.5 5</intersection>
<intersection>-14 3</intersection>
<intersection>15 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,21,23,21</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,15,18.5,15</points>
<connection>
<GID>58</GID>
<name>Q</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>18.5,-14,221.5,-14</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>18.5,-23.5,37.5,-23.5</points>
<intersection>18.5 0</intersection>
<intersection>37.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>37.5,-56,37.5,-23.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-23.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>18.5,-29.5,24.5,-29.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,5.5,14.5,11</points>
<intersection>5.5 3</intersection>
<intersection>11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,11,14.5,11</points>
<connection>
<GID>58</GID>
<name>nQ</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14.5,5.5,22,5.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,13.5,33,23</points>
<intersection>13.5 1</intersection>
<intersection>22 2</intersection>
<intersection>23 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,13.5,37,13.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,22,33,22</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,23,64,23</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,2.5,33.5,11.5</points>
<intersection>2.5 2</intersection>
<intersection>4.5 3</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,11.5,37,11.5</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,2.5,66.5,2.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,4.5,33.5,4.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-55.5,63,21</points>
<intersection>-55.5 9</intersection>
<intersection>-29 5</intersection>
<intersection>-13 3</intersection>
<intersection>14.5 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,21,64,21</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,14.5,63,14.5</points>
<connection>
<GID>60</GID>
<name>Q</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>63,-13,221.5,-13</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-29,67.5,-29</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>50,-55.5,63,-55.5</points>
<intersection>50 10</intersection>
<intersection>63 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>50,-57,50,-55.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-55.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-44.5,47,-29.5</points>
<intersection>-44.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-29.5,47,-29.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-44.5,241,-44.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,21.5,71.5,22</points>
<intersection>21.5 2</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,22,71.5,22</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,21.5,93.5,21.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection>
<intersection>73.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>73.5,14.5,73.5,21.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>21.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,4.5,64.5,10.5</points>
<intersection>4.5 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,10.5,64.5,10.5</points>
<connection>
<GID>60</GID>
<name>nQ</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,4.5,66.5,4.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,1,73,12.5</points>
<intersection>1 3</intersection>
<intersection>3.5 1</intersection>
<intersection>12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,3.5,73,3.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,12.5,73.5,12.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>73,1,96,1</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-56,90,41.5</points>
<intersection>-56 13</intersection>
<intersection>-29 9</intersection>
<intersection>-12 2</intersection>
<intersection>15 1</intersection>
<intersection>19.5 5</intersection>
<intersection>41.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,15,90,15</points>
<connection>
<GID>63</GID>
<name>Q</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90,-12,221.5,-12</points>
<connection>
<GID>109</GID>
<name>IN_2</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>90,19.5,93.5,19.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>90,41.5,223.5,41.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>90,-29,97,-29</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>90,-56,114,-56</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,20.5,120,20.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,14,102,20.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,1,102,12</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,1,121.5,1</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,3,91.5,11</points>
<intersection>3 2</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,11,91.5,11</points>
<connection>
<GID>63</GID>
<name>nQ</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,3,96,3</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-29,118,39.5</points>
<connection>
<GID>65</GID>
<name>Q</name></connection>
<intersection>-29 10</intersection>
<intersection>-11 2</intersection>
<intersection>18.5 6</intersection>
<intersection>39.5 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>118,-11,221.5,-11</points>
<connection>
<GID>109</GID>
<name>IN_3</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>118,18.5,120,18.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118,39.5,223.5,39.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>118,-29,125.5,-29</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection>
<intersection>121 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>121,-56,121,-29</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-29 10</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,3,119,10.5</points>
<intersection>3 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,10.5,119,10.5</points>
<connection>
<GID>65</GID>
<name>nQ</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,3,121.5,3</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,13.5,129,21.5</points>
<intersection>13.5 2</intersection>
<intersection>19.5 1</intersection>
<intersection>21.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,19.5,129,19.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129,13.5,131,13.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129,21.5,167,21.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,2,129.5,11.5</points>
<intersection>2 1</intersection>
<intersection>11.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,2,167.5,2</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>129.5,11.5,131,11.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-55.5,161.5,37.5</points>
<intersection>-55.5 14</intersection>
<intersection>-29 9</intersection>
<intersection>-10 3</intersection>
<intersection>12.5 1</intersection>
<intersection>19.5 10</intersection>
<intersection>37.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,12.5,161.5,12.5</points>
<connection>
<GID>67</GID>
<name>Q</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>161.5,-10,221.5,-10</points>
<connection>
<GID>109</GID>
<name>IN_4</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>161.5,37.5,223.5,37.5</points>
<connection>
<GID>51</GID>
<name>IN_2</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>161.5,-29,171.5,-29</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>161.5,19.5,167,19.5</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>161.5,-55.5,178.5,-55.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,4,159,8.5</points>
<intersection>4 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,8.5,159,8.5</points>
<connection>
<GID>67</GID>
<name>nQ</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>159,4,167.5,4</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,13,174,20.5</points>
<intersection>13 2</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,20.5,174,20.5</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,13,175,13</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,3,174,11</points>
<intersection>3 1</intersection>
<intersection>11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,3,174,3</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,11,175,11</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-6.5,199,-6.5</points>
<intersection>-19 16</intersection>
<intersection>-1.5 13</intersection>
<intersection>55.5 12</intersection>
<intersection>81 6</intersection>
<intersection>109 7</intersection>
<intersection>147 11</intersection>
<intersection>199 28</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>81,-6.5,81,13</points>
<intersection>-6.5 1</intersection>
<intersection>13 19</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>109,-6.5,109,12.5</points>
<intersection>-6.5 1</intersection>
<intersection>12.5 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>147,-6.5,147,10.5</points>
<intersection>-6.5 1</intersection>
<intersection>10.5 18</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>55.5,-6.5,55.5,12.5</points>
<intersection>-6.5 1</intersection>
<intersection>12.5 22</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-1.5,-6.5,-1.5,13</points>
<intersection>-6.5 1</intersection>
<intersection>13 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>109,12.5,112,12.5</points>
<connection>
<GID>65</GID>
<name>clock</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-1.5,13,6.5,13</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>-1.5 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-19,-36,-19,-6.5</points>
<intersection>-36 17</intersection>
<intersection>-7 37</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-19,-36,219.5,-36</points>
<intersection>-19 16</intersection>
<intersection>24.5 34</intersection>
<intersection>67.5 25</intersection>
<intersection>97 26</intersection>
<intersection>125.5 24</intersection>
<intersection>170.5 23</intersection>
<intersection>219.5 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>147,10.5,150.5,10.5</points>
<connection>
<GID>67</GID>
<name>clock</name></connection>
<intersection>147 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>81,13,82,13</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>81 6</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>55.5,12.5,56,12.5</points>
<connection>
<GID>60</GID>
<name>clock</name></connection>
<intersection>55.5 12</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>170.5,-36,170.5,-32</points>
<intersection>-36 17</intersection>
<intersection>-32 36</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>125.5,-36,125.5,-32</points>
<connection>
<GID>86</GID>
<name>clock</name></connection>
<intersection>-36 17</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>67.5,-36,67.5,-32</points>
<connection>
<GID>61</GID>
<name>clock</name></connection>
<intersection>-36 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>97,-36,97,-32</points>
<connection>
<GID>73</GID>
<name>clock</name></connection>
<intersection>-36 17</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>199,-6.5,199,10</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>-6.5 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>24.5,-36,24.5,-32.5</points>
<connection>
<GID>57</GID>
<name>clock</name></connection>
<intersection>-36 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>219.5,-36,219.5,-32.5</points>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<intersection>-36 17</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>170.5,-32,171.5,-32</points>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<intersection>170.5 23</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-60,-7,-19,-7</points>
<connection>
<GID>501</GID>
<name>OUT</name></connection>
<intersection>-57.5 38</intersection>
<intersection>-19 16</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>-57.5,-7,-57.5,3.5</points>
<intersection>-7 37</intersection>
<intersection>3.5 39</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-57.5,3.5,-57,3.5</points>
<connection>
<GID>496</GID>
<name>clock</name></connection>
<intersection>-57.5 38</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-55,214,35.5</points>
<intersection>-55 9</intersection>
<intersection>-29.5 13</intersection>
<intersection>-9 2</intersection>
<intersection>12 11</intersection>
<intersection>35.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>214,-9,221.5,-9</points>
<connection>
<GID>109</GID>
<name>IN_5</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>214,35.5,223.5,35.5</points>
<connection>
<GID>51</GID>
<name>IN_3</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>184,-55,214,-55</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>205,12,214,12</points>
<connection>
<GID>69</GID>
<name>Q</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>214,-29.5,219.5,-29.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>214 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-43.5,241,-43.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>75 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-43.5,75,-29</points>
<intersection>-43.5 1</intersection>
<intersection>-29 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-29,75,-29</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>75 3</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-42.5,241,-42.5</points>
<connection>
<GID>111</GID>
<name>IN_2</name></connection>
<intersection>104.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>104.5,-42.5,104.5,-29</points>
<intersection>-42.5 1</intersection>
<intersection>-29 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>103,-29,104.5,-29</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>104.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-41.5,241,-41.5</points>
<connection>
<GID>111</GID>
<name>IN_3</name></connection>
<intersection>131.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-41.5,131.5,-29</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-40.5,184,-29</points>
<intersection>-40.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177.5,-29,184,-29</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184,-40.5,241,-40.5</points>
<connection>
<GID>111</GID>
<name>IN_4</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>232.5,-39.5,241,-39.5</points>
<connection>
<GID>111</GID>
<name>IN_5</name></connection>
<intersection>232.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>232.5,-39.5,232.5,-29.5</points>
<intersection>-39.5 1</intersection>
<intersection>-29.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>225.5,-29.5,232.5,-29.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>232.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,15,3.5,27.5</points>
<intersection>15 8</intersection>
<intersection>27.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-5,27.5,3.5,27.5</points>
<intersection>-5 9</intersection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>3.5,15,6.5,15</points>
<connection>
<GID>58</GID>
<name>J</name></connection>
<intersection>3.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-5,27,-5,39</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>27.5 6</intersection>
<intersection>39 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-46,39,-5,39</points>
<intersection>-46 14</intersection>
<intersection>-5 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-46,35.5,-46,39</points>
<intersection>35.5 15</intersection>
<intersection>39 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-56.5,35.5,-46,35.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>-46 14</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-11.5,34.5,186.5,34.5</points>
<intersection>-11.5 7</intersection>
<intersection>44 6</intersection>
<intersection>80.5 10</intersection>
<intersection>109 12</intersection>
<intersection>139 14</intersection>
<intersection>186.5 16</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>44,29.5,44,34.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>34.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-11.5,27.5,-11.5,34.5</points>
<intersection>27.5 20</intersection>
<intersection>34.5 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>80.5,30,80.5,34.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>34.5 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>109,29.5,109,34.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>34.5 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>139,29.5,139,34.5</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>34.5 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>186.5,31.5,186.5,34.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>34.5 4</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-42,27.5,-7,27.5</points>
<intersection>-42 23</intersection>
<intersection>-11.5 7</intersection>
<intersection>-7 26</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-42,-108,-42,27.5</points>
<intersection>-108 24</intersection>
<intersection>27.5 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-42,-108,22,-108</points>
<intersection>-42 23</intersection>
<intersection>22 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>22,-108,22,-107</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-108 24</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-7,27,-7,27.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>27.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,11,-6,21</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,11,6.5,11</points>
<connection>
<GID>58</GID>
<name>K</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-66.5,41.5,-57.5,41.5</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,41.5,-55.5,42.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>42.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-49.5,42.5,-49.5,44</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,42.5,-49.5,42.5</points>
<intersection>-55.5 0</intersection>
<intersection>-49.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-79,42.5,-67.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-67.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>37.5,-67.5,37.5,-62</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-67.5,42.5,-67.5</points>
<intersection>37.5 1</intersection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-79,44.5,-67.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-67.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-67.5,50,-63</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-67.5,50,-67.5</points>
<intersection>44.5 0</intersection>
<intersection>50 1</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-101,21,-88.5</points>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>43.5,-88.5,43.5,-85</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>21,-88.5,43.5,-88.5</points>
<intersection>21 0</intersection>
<intersection>43.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-65.5,118.5,-63.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>121,-63.5,121,-62</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>118.5,-63.5,121,-63.5</points>
<intersection>118.5 0</intersection>
<intersection>121 1</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-65.5,116.5,-63.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>114,-63.5,114,-62</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>114,-63.5,116.5,-63.5</points>
<intersection>114 1</intersection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-101,23,-90.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>117.5,-90.5,117.5,-71.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23,-90.5,117.5,-90.5</points>
<intersection>23 0</intersection>
<intersection>117.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-64,181.5,-62.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>184,-62.5,184,-61</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-62.5,184,-62.5</points>
<intersection>181.5 0</intersection>
<intersection>184 1</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-64,179.5,-62.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>178.5,-62.5,178.5,-61.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-62.5,179.5,-62.5</points>
<intersection>178.5 1</intersection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-101,25,-93</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>180.5,-93,180.5,-70</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-93,180.5,-93</points>
<intersection>25 0</intersection>
<intersection>180.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,12.5,53.5,30</points>
<intersection>12.5 2</intersection>
<intersection>14.5 1</intersection>
<intersection>30 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,14.5,56,14.5</points>
<connection>
<GID>60</GID>
<name>J</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,12.5,53.5,12.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46,30,53.5,30</points>
<intersection>46 4</intersection>
<intersection>53.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46,29.5,46,30</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>30 3</intersection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,10.5,45,23.5</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,10.5,56,10.5</points>
<connection>
<GID>60</GID>
<name>K</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,15,81.5,24</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,15,82,15</points>
<connection>
<GID>63</GID>
<name>J</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,22.5,89,30</points>
<intersection>22.5 1</intersection>
<intersection>30 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,22.5,89,22.5</points>
<intersection>79.5 4</intersection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>82.5,30,89,30</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>79.5,11,79.5,22.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>11 6</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>79.5,11,82,11</points>
<connection>
<GID>63</GID>
<name>K</name></connection>
<intersection>79.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,22,114.5,22</points>
<intersection>108 3</intersection>
<intersection>114.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,13,108,22</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>14.5 7</intersection>
<intersection>22 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>114.5,22,114.5,29.5</points>
<intersection>22 1</intersection>
<intersection>29.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>111,29.5,114.5,29.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>114.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>108,14.5,112,14.5</points>
<connection>
<GID>65</GID>
<name>J</name></connection>
<intersection>108 3</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,10.5,110,23.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,10.5,112,10.5</points>
<connection>
<GID>65</GID>
<name>K</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,12.5,150.5,12.5</points>
<connection>
<GID>67</GID>
<name>J</name></connection>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>148 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>148,12.5,148,30.5</points>
<intersection>12.5 1</intersection>
<intersection>30.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>141,30.5,148,30.5</points>
<intersection>141 6</intersection>
<intersection>148 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>141,29.5,141,30.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>30.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,8.5,140,23.5</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,8.5,150.5,8.5</points>
<connection>
<GID>67</GID>
<name>K</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181,12,199,12</points>
<connection>
<GID>69</GID>
<name>J</name></connection>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>193.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>193.5,12,193.5,33</points>
<intersection>12 1</intersection>
<intersection>33 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>188.5,33,193.5,33</points>
<intersection>188.5 15</intersection>
<intersection>193.5 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>188.5,31.5,188.5,33</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>33 8</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,8,187.5,25.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,8,199,8</points>
<connection>
<GID>69</GID>
<name>K</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-767.429,20.8773,295.904,-504.708</PageViewport>
<gate>
<ID>788</ID>
<type>AE_DFF_LOW</type>
<position>-97,-426.5</position>
<input>
<ID>IN_0</ID>805 </input>
<output>
<ID>OUT_0</ID>811 </output>
<input>
<ID>clock</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>789</ID>
<type>AE_DFF_LOW</type>
<position>-81,-427</position>
<input>
<ID>IN_0</ID>806 </input>
<output>
<ID>OUT_0</ID>812 </output>
<input>
<ID>clock</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>790</ID>
<type>AE_DFF_LOW</type>
<position>-67.5,-427</position>
<input>
<ID>IN_0</ID>807 </input>
<output>
<ID>OUT_0</ID>813 </output>
<input>
<ID>clock</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>791</ID>
<type>AE_DFF_LOW</type>
<position>-52.5,-427</position>
<input>
<ID>IN_0</ID>808 </input>
<output>
<ID>OUT_0</ID>814 </output>
<input>
<ID>clock</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>792</ID>
<type>AE_DFF_LOW</type>
<position>-42,-427</position>
<input>
<ID>IN_0</ID>809 </input>
<output>
<ID>OUT_0</ID>815 </output>
<input>
<ID>clock</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>793</ID>
<type>AE_DFF_LOW</type>
<position>-29,-427</position>
<input>
<ID>IN_0</ID>810 </input>
<output>
<ID>OUT_0</ID>816 </output>
<input>
<ID>clock</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>794</ID>
<type>AE_SMALL_INVERTER</type>
<position>-90,-434.5</position>
<input>
<ID>IN_0</ID>811 </input>
<output>
<ID>OUT_0</ID>817 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>795</ID>
<type>AE_SMALL_INVERTER</type>
<position>-75,-434.5</position>
<input>
<ID>IN_0</ID>812 </input>
<output>
<ID>OUT_0</ID>818 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>796</ID>
<type>AE_SMALL_INVERTER</type>
<position>-60,-434.5</position>
<input>
<ID>IN_0</ID>813 </input>
<output>
<ID>OUT_0</ID>819 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>797</ID>
<type>AE_SMALL_INVERTER</type>
<position>-48.5,-434</position>
<input>
<ID>IN_0</ID>814 </input>
<output>
<ID>OUT_0</ID>820 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>798</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35.5,-434.5</position>
<input>
<ID>IN_0</ID>815 </input>
<output>
<ID>OUT_0</ID>821 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>799</ID>
<type>AE_SMALL_INVERTER</type>
<position>-22.5,-434</position>
<input>
<ID>IN_0</ID>816 </input>
<output>
<ID>OUT_0</ID>822 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_AND4</type>
<position>-72,-451</position>
<input>
<ID>IN_0</ID>820 </input>
<input>
<ID>IN_1</ID>819 </input>
<input>
<ID>IN_2</ID>818 </input>
<input>
<ID>IN_3</ID>817 </input>
<output>
<ID>OUT</ID>823 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>801</ID>
<type>AA_AND2</type>
<position>-35.5,-450</position>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>821 </input>
<output>
<ID>OUT</ID>824 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>802</ID>
<type>AA_AND2</type>
<position>-56.5,-463</position>
<input>
<ID>IN_0</ID>824 </input>
<input>
<ID>IN_1</ID>823 </input>
<output>
<ID>OUT</ID>827 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>803</ID>
<type>AI_XOR2</type>
<position>-581,-14.5</position>
<input>
<ID>IN_0</ID>827 </input>
<input>
<ID>IN_1</ID>825 </input>
<output>
<ID>OUT</ID>826 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>804</ID>
<type>AA_LABEL</type>
<position>-507,-208.5</position>
<gparam>LABEL_TEXT Default Power</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>805</ID>
<type>AE_DFF_LOW</type>
<position>-595.5,-200</position>
<input>
<ID>IN_0</ID>829 </input>
<output>
<ID>OUTINV_0</ID>831 </output>
<output>
<ID>OUT_0</ID>887 </output>
<input>
<ID>clear</ID>835 </input>
<input>
<ID>clock</ID>830 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>806</ID>
<type>BB_CLOCK</type>
<position>-610.5,-203.5</position>
<output>
<ID>CLK</ID>830 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>807</ID>
<type>AA_LABEL</type>
<position>-478,-337</position>
<gparam>LABEL_TEXT Checking condition for 60</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>808</ID>
<type>AA_TOGGLE</type>
<position>-608.5,-198</position>
<output>
<ID>OUT_0</ID>829 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>809</ID>
<type>AA_LABEL</type>
<position>-276.5,-256</position>
<gparam>LABEL_TEXT Problematic Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>810</ID>
<type>BA_NAND4</type>
<position>-299.5,-201</position>
<input>
<ID>IN_0</ID>846 </input>
<input>
<ID>IN_1</ID>850 </input>
<input>
<ID>IN_2</ID>854 </input>
<input>
<ID>IN_3</ID>859 </input>
<output>
<ID>OUT</ID>836 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>811</ID>
<type>AE_DFF_LOW</type>
<position>-498.5,-271</position>
<input>
<ID>IN_0</ID>837 </input>
<output>
<ID>OUT_0</ID>842 </output>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>812</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-516.5,-226.5</position>
<input>
<ID>J</ID>865 </input>
<input>
<ID>K</ID>867 </input>
<output>
<ID>Q</ID>837 </output>
<input>
<ID>clear</ID>836 </input>
<input>
<ID>clock</ID>858 </input>
<output>
<ID>nQ</ID>838 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>813</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-467,-227</position>
<input>
<ID>J</ID>877 </input>
<input>
<ID>K</ID>878 </input>
<output>
<ID>Q</ID>841 </output>
<input>
<ID>clear</ID>836 </input>
<input>
<ID>clock</ID>858 </input>
<output>
<ID>nQ</ID>844 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>814</ID>
<type>AE_DFF_LOW</type>
<position>-455.5,-270.5</position>
<input>
<ID>IN_0</ID>841 </input>
<output>
<ID>OUT_0</ID>860 </output>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>815</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-441,-226.5</position>
<input>
<ID>J</ID>879 </input>
<input>
<ID>K</ID>880 </input>
<output>
<ID>Q</ID>846 </output>
<input>
<ID>clear</ID>836 </input>
<input>
<ID>clock</ID>858 </input>
<output>
<ID>nQ</ID>849 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>816</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-411,-227</position>
<input>
<ID>J</ID>881 </input>
<input>
<ID>K</ID>882 </input>
<output>
<ID>Q</ID>850 </output>
<input>
<ID>clear</ID>836 </input>
<input>
<ID>clock</ID>858 </input>
<output>
<ID>nQ</ID>851 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>817</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-372.5,-229</position>
<input>
<ID>J</ID>883 </input>
<input>
<ID>K</ID>884 </input>
<output>
<ID>Q</ID>854 </output>
<input>
<ID>clear</ID>836 </input>
<input>
<ID>clock</ID>858 </input>
<output>
<ID>nQ</ID>855 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>818</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-324,-229.5</position>
<input>
<ID>J</ID>885 </input>
<input>
<ID>K</ID>886 </input>
<output>
<ID>Q</ID>859 </output>
<input>
<ID>clear</ID>836 </input>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>819</ID>
<type>AE_DFF_LOW</type>
<position>-426,-270.5</position>
<input>
<ID>IN_0</ID>846 </input>
<output>
<ID>OUT_0</ID>861 </output>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>820</ID>
<type>AA_AND2</type>
<position>-500,-217.5</position>
<input>
<ID>IN_0</ID>893 </input>
<input>
<ID>IN_1</ID>837 </input>
<output>
<ID>OUT</ID>839 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>821</ID>
<type>AA_AND2</type>
<position>-501,-235</position>
<input>
<ID>IN_0</ID>838 </input>
<input>
<ID>IN_1</ID>894 </input>
<output>
<ID>OUT</ID>840 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>822</ID>
<type>AA_AND2</type>
<position>-459,-217.5</position>
<input>
<ID>IN_0</ID>839 </input>
<input>
<ID>IN_1</ID>841 </input>
<output>
<ID>OUT</ID>843 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>823</ID>
<type>AA_AND2</type>
<position>-456.5,-236</position>
<input>
<ID>IN_0</ID>844 </input>
<input>
<ID>IN_1</ID>840 </input>
<output>
<ID>OUT</ID>845 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>824</ID>
<type>AA_AND2</type>
<position>-429.5,-219</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>846 </input>
<output>
<ID>OUT</ID>847 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>825</ID>
<type>AA_AND2</type>
<position>-427,-237.5</position>
<input>
<ID>IN_0</ID>849 </input>
<input>
<ID>IN_1</ID>845 </input>
<output>
<ID>OUT</ID>848 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>826</ID>
<type>AA_AND2</type>
<position>-403,-220</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>850 </input>
<output>
<ID>OUT</ID>852 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>827</ID>
<type>AA_AND2</type>
<position>-401.5,-237.5</position>
<input>
<ID>IN_0</ID>851 </input>
<input>
<ID>IN_1</ID>848 </input>
<output>
<ID>OUT</ID>853 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>828</ID>
<type>AA_AND2</type>
<position>-356,-219</position>
<input>
<ID>IN_0</ID>852 </input>
<input>
<ID>IN_1</ID>854 </input>
<output>
<ID>OUT</ID>856 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>829</ID>
<type>AA_AND2</type>
<position>-355.5,-236.5</position>
<input>
<ID>IN_0</ID>855 </input>
<input>
<ID>IN_1</ID>853 </input>
<output>
<ID>OUT</ID>857 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>830</ID>
<type>AE_DFF_LOW</type>
<position>-397.5,-270.5</position>
<input>
<ID>IN_0</ID>850 </input>
<output>
<ID>OUT_0</ID>862 </output>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>831</ID>
<type>AE_OR2</type>
<position>-486,-227</position>
<input>
<ID>IN_0</ID>839 </input>
<input>
<ID>IN_1</ID>840 </input>
<output>
<ID>OUT</ID>877 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>832</ID>
<type>AE_DFF_LOW</type>
<position>-351.5,-270.5</position>
<input>
<ID>IN_0</ID>854 </input>
<output>
<ID>OUT_0</ID>863 </output>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>833</ID>
<type>AE_OR2</type>
<position>-449.5,-226</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>845 </input>
<output>
<ID>OUT</ID>880 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>834</ID>
<type>AE_OR2</type>
<position>-421,-226.5</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>848 </input>
<output>
<ID>OUT</ID>881 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>835</ID>
<type>AE_OR2</type>
<position>-392,-227</position>
<input>
<ID>IN_0</ID>852 </input>
<input>
<ID>IN_1</ID>853 </input>
<output>
<ID>OUT</ID>883 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>836</ID>
<type>AE_OR2</type>
<position>-348,-227.5</position>
<input>
<ID>IN_0</ID>856 </input>
<input>
<ID>IN_1</ID>857 </input>
<output>
<ID>OUT</ID>885 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>837</ID>
<type>AE_DFF_LOW</type>
<position>-303.5,-271</position>
<input>
<ID>IN_0</ID>859 </input>
<output>
<ID>OUT_0</ID>864 </output>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>838</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-299.5,-250.5</position>
<input>
<ID>IN_0</ID>837 </input>
<input>
<ID>IN_1</ID>841 </input>
<input>
<ID>IN_2</ID>846 </input>
<input>
<ID>IN_3</ID>850 </input>
<input>
<ID>IN_4</ID>854 </input>
<input>
<ID>IN_5</ID>859 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>839</ID>
<type>AE_DFF_LOW</type>
<position>-580,-235</position>
<input>
<ID>IN_0</ID>892 </input>
<output>
<ID>OUTINV_0</ID>894 </output>
<output>
<ID>OUT_0</ID>893 </output>
<input>
<ID>clear</ID>835 </input>
<input>
<ID>clock</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>840</ID>
<type>CC_PULSE</type>
<position>-626,-229.5</position>
<output>
<ID>OUT_0</ID>890 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>841</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-280,-281</position>
<input>
<ID>IN_0</ID>842 </input>
<input>
<ID>IN_1</ID>860 </input>
<input>
<ID>IN_2</ID>861 </input>
<input>
<ID>IN_3</ID>862 </input>
<input>
<ID>IN_4</ID>863 </input>
<input>
<ID>IN_5</ID>864 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 21</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>842</ID>
<type>CC_PULSE</type>
<position>-626,-247.5</position>
<output>
<ID>OUT_0</ID>889 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>843</ID>
<type>EE_VDD</type>
<position>-575.5,-194.5</position>
<output>
<ID>OUT_0</ID>888 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>844</ID>
<type>AE_OR2</type>
<position>-589,-246.5</position>
<input>
<ID>IN_0</ID>890 </input>
<input>
<ID>IN_1</ID>889 </input>
<output>
<ID>OUT</ID>858 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>845</ID>
<type>AE_SMALL_INVERTER</type>
<position>-606.5,-230</position>
<input>
<ID>IN_0</ID>890 </input>
<output>
<ID>OUT_0</ID>891 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>846</ID>
<type>AA_AND2</type>
<position>-482.5,-321.5</position>
<input>
<ID>IN_0</ID>869 </input>
<input>
<ID>IN_1</ID>868 </input>
<output>
<ID>OUT</ID>870 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>847</ID>
<type>AI_XOR2</type>
<position>-592,-234</position>
<input>
<ID>IN_0</ID>889 </input>
<input>
<ID>IN_1</ID>891 </input>
<output>
<ID>OUT</ID>892 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>848</ID>
<type>AA_LABEL</type>
<position>-622,-223.5</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>849</ID>
<type>AA_AND2</type>
<position>-408.5,-308</position>
<input>
<ID>IN_0</ID>871 </input>
<input>
<ID>IN_1</ID>872 </input>
<output>
<ID>OUT</ID>873 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>850</ID>
<type>AA_LABEL</type>
<position>-623,-252.5</position>
<gparam>LABEL_TEXT Decrement</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>851</ID>
<type>AA_AND2</type>
<position>-345.5,-306.5</position>
<input>
<ID>IN_0</ID>874 </input>
<input>
<ID>IN_1</ID>875 </input>
<output>
<ID>OUT</ID>876 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>852</ID>
<type>AI_XOR2</type>
<position>-532,-215.5</position>
<input>
<ID>IN_0</ID>865 </input>
<input>
<ID>IN_1</ID>866 </input>
<output>
<ID>OUT</ID>867 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>853</ID>
<type>AI_XOR2</type>
<position>-481,-213</position>
<input>
<ID>IN_0</ID>877 </input>
<input>
<ID>IN_1</ID>866 </input>
<output>
<ID>OUT</ID>878 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>854</ID>
<type>AI_XOR2</type>
<position>-444.5,-212.5</position>
<input>
<ID>IN_0</ID>880 </input>
<input>
<ID>IN_1</ID>866 </input>
<output>
<ID>OUT</ID>879 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>855</ID>
<type>AI_XOR2</type>
<position>-416,-213</position>
<input>
<ID>IN_0</ID>881 </input>
<input>
<ID>IN_1</ID>866 </input>
<output>
<ID>OUT</ID>882 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>856</ID>
<type>AI_XOR2</type>
<position>-386,-213</position>
<input>
<ID>IN_0</ID>883 </input>
<input>
<ID>IN_1</ID>866 </input>
<output>
<ID>OUT</ID>884 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>857</ID>
<type>AI_XOR2</type>
<position>-338.5,-211</position>
<input>
<ID>IN_0</ID>885 </input>
<input>
<ID>IN_1</ID>866 </input>
<output>
<ID>OUT</ID>886 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>858</ID>
<type>AA_AND4</type>
<position>-504,-343.5</position>
<input>
<ID>IN_0</ID>876 </input>
<input>
<ID>IN_1</ID>873 </input>
<input>
<ID>IN_2</ID>870 </input>
<input>
<ID>IN_3</ID>894 </input>
<output>
<ID>OUT</ID>866 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>859</ID>
<type>AA_INVERTER</type>
<position>-488.5,-298.5</position>
<input>
<ID>IN_0</ID>837 </input>
<output>
<ID>OUT_0</ID>868 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>860</ID>
<type>AA_INVERTER</type>
<position>-476,-299.5</position>
<input>
<ID>IN_0</ID>841 </input>
<output>
<ID>OUT_0</ID>869 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>861</ID>
<type>AA_INVERTER</type>
<position>-412,-298.5</position>
<input>
<ID>IN_0</ID>846 </input>
<output>
<ID>OUT_0</ID>872 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>862</ID>
<type>AA_INVERTER</type>
<position>-405,-298.5</position>
<input>
<ID>IN_0</ID>850 </input>
<output>
<ID>OUT_0</ID>871 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>863</ID>
<type>AA_INVERTER</type>
<position>-347.5,-298</position>
<input>
<ID>IN_0</ID>854 </input>
<output>
<ID>OUT_0</ID>875 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>864</ID>
<type>AA_INVERTER</type>
<position>-342,-297.5</position>
<input>
<ID>IN_0</ID>859 </input>
<output>
<ID>OUT_0</ID>874 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>865</ID>
<type>AA_LABEL</type>
<position>-280,-291</position>
<gparam>LABEL_TEXT Actual Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>866</ID>
<type>AA_LABEL</type>
<position>-558.5,-254</position>
<gparam>LABEL_TEXT Clock input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>867</ID>
<type>AA_AND2</type>
<position>-582.5,-201</position>
<input>
<ID>IN_0</ID>888 </input>
<input>
<ID>IN_1</ID>887 </input>
<output>
<ID>OUT</ID>865 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>868</ID>
<type>AA_LABEL</type>
<position>-453.5,-191.5</position>
<gparam>LABEL_TEXT Setting Mode</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>869</ID>
<type>AA_LABEL</type>
<position>-588.5,-188</position>
<gparam>LABEL_TEXT On/Off- Settings/Cycle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>870</ID>
<type>AA_LABEL</type>
<position>-559,-222.5</position>
<gparam>LABEL_TEXT Direction</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>871</ID>
<type>AA_INVERTER</type>
<position>-412,-75</position>
<input>
<ID>IN_0</ID>945 </input>
<output>
<ID>OUT_0</ID>898 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>872</ID>
<type>AA_LABEL</type>
<position>-602,0.5</position>
<gparam>LABEL_TEXT Water Button</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>873</ID>
<type>AA_LABEL</type>
<position>-451.5,-40.5</position>
<gparam>LABEL_TEXT Buffer Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>874</ID>
<type>AA_LABEL</type>
<position>-509.5,11</position>
<gparam>LABEL_TEXT Seconds Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>875</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-322.5,-102</position>
<input>
<ID>J</ID>898 </input>
<input>
<ID>K</ID>906 </input>
<output>
<ID>Q</ID>896 </output>
<input>
<ID>clock</ID>917 </input>
<output>
<ID>nQ</ID>902 </output>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>876</ID>
<type>AA_LABEL</type>
<position>-453,-62</position>
<gparam>LABEL_TEXT Actual Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>877</ID>
<type>AA_LABEL</type>
<position>-379,-80.5</position>
<gparam>LABEL_TEXT Minutes Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>878</ID>
<type>AA_LABEL</type>
<position>-316,-116</position>
<gparam>LABEL_TEXT Buffer Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>879</ID>
<type>AI_XOR2</type>
<position>-437,-16</position>
<input>
<ID>IN_0</ID>902 </input>
<input>
<ID>IN_1</ID>904 </input>
<output>
<ID>OUT</ID>910 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>880</ID>
<type>AA_LABEL</type>
<position>-432.5,-6</position>
<gparam>LABEL_TEXT Both on seconds counter stop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>881</ID>
<type>AA_LABEL</type>
<position>-306.5,-145</position>
<gparam>LABEL_TEXT Actual Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>882</ID>
<type>AI_XOR2</type>
<position>-338,-104</position>
<input>
<ID>IN_0</ID>911 </input>
<input>
<ID>IN_1</ID>896 </input>
<output>
<ID>OUT</ID>899 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>883</ID>
<type>AA_INVERTER</type>
<position>-329,-87</position>
<input>
<ID>IN_0</ID>905 </input>
<output>
<ID>OUT_0</ID>906 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>884</ID>
<type>AA_AND2</type>
<position>-575.5,-39.5</position>
<input>
<ID>IN_0</ID>945 </input>
<input>
<ID>IN_1</ID>895 </input>
<output>
<ID>OUT</ID>917 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>885</ID>
<type>AA_LABEL</type>
<position>-586.5,-113.5</position>
<gparam>LABEL_TEXT Abort</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>886</ID>
<type>AE_OR2</type>
<position>-522,-95.5</position>
<input>
<ID>IN_0</ID>928 </input>
<input>
<ID>IN_1</ID>927 </input>
<output>
<ID>OUT</ID>900 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>887</ID>
<type>AA_TOGGLE</type>
<position>-586,-108.5</position>
<output>
<ID>OUT_0</ID>911 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>888</ID>
<type>AE_OR4</type>
<position>-554,-87</position>
<input>
<ID>IN_0</ID>926 </input>
<input>
<ID>IN_1</ID>925 </input>
<input>
<ID>IN_2</ID>924 </input>
<input>
<ID>IN_3</ID>923 </input>
<output>
<ID>OUT</ID>897 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>889</ID>
<type>AE_OR2</type>
<position>-568,-92.5</position>
<input>
<ID>IN_0</ID>900 </input>
<input>
<ID>IN_1</ID>897 </input>
<output>
<ID>OUT</ID>907 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>890</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-563,-27</position>
<input>
<ID>J</ID>945 </input>
<input>
<ID>K</ID>945 </input>
<output>
<ID>Q</ID>916 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>891</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-549.5,-27</position>
<input>
<ID>J</ID>916 </input>
<input>
<ID>K</ID>916 </input>
<output>
<ID>Q</ID>918 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>892</ID>
<type>AA_AND2</type>
<position>-574.5,-83</position>
<input>
<ID>IN_0</ID>899 </input>
<input>
<ID>IN_1</ID>945 </input>
<output>
<ID>OUT</ID>901 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>893</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-533.5,-27</position>
<input>
<ID>J</ID>912 </input>
<input>
<ID>K</ID>912 </input>
<output>
<ID>Q</ID>920 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>894</ID>
<type>AE_OR2</type>
<position>-593,-80</position>
<input>
<ID>IN_0</ID>908 </input>
<input>
<ID>IN_1</ID>901 </input>
<output>
<ID>OUT</ID>909 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>895</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-517.5,-27.5</position>
<input>
<ID>J</ID>913 </input>
<input>
<ID>K</ID>913 </input>
<output>
<ID>Q</ID>919 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>896</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-501.5,-28</position>
<input>
<ID>J</ID>914 </input>
<input>
<ID>K</ID>914 </input>
<output>
<ID>Q</ID>921 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>897</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-484.5,-28</position>
<input>
<ID>J</ID>915 </input>
<input>
<ID>K</ID>915 </input>
<output>
<ID>Q</ID>922 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>898</ID>
<type>AI_XOR2</type>
<position>-452,-25</position>
<input>
<ID>IN_0</ID>911 </input>
<input>
<ID>IN_1</ID>910 </input>
<output>
<ID>OUT</ID>903 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>899</ID>
<type>AA_TOGGLE</type>
<position>-593.5,-7</position>
<output>
<ID>OUT_0</ID>825 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>900</ID>
<type>AA_LABEL</type>
<position>-606.5,-73</position>
<gparam>LABEL_TEXT Water On/Off</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>901</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-434.5,-100</position>
<input>
<ID>J</ID>945 </input>
<input>
<ID>K</ID>945 </input>
<output>
<ID>Q</ID>933 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>902</ID>
<type>AA_AND2</type>
<position>-585.5,-91.5</position>
<input>
<ID>IN_0</ID>907 </input>
<input>
<ID>IN_1</ID>945 </input>
<output>
<ID>OUT</ID>908 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>903</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-421,-100</position>
<input>
<ID>J</ID>933 </input>
<input>
<ID>K</ID>933 </input>
<output>
<ID>Q</ID>934 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>904</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-467,-41.5</position>
<input>
<ID>IN_0</ID>916 </input>
<input>
<ID>IN_1</ID>918 </input>
<input>
<ID>IN_2</ID>920 </input>
<input>
<ID>IN_3</ID>919 </input>
<input>
<ID>IN_4</ID>921 </input>
<input>
<ID>IN_5</ID>922 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>905</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-405,-100</position>
<input>
<ID>J</ID>929 </input>
<input>
<ID>K</ID>929 </input>
<output>
<ID>Q</ID>936 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>906</ID>
<type>GA_LED</type>
<position>-605,-80</position>
<input>
<ID>N_in1</ID>909 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>907</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-389,-100.5</position>
<input>
<ID>J</ID>930 </input>
<input>
<ID>K</ID>930 </input>
<output>
<ID>Q</ID>935 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>908</ID>
<type>AA_LABEL</type>
<position>-554.5,-98</position>
<gparam>LABEL_TEXT Output of Flip-flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>909</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-373,-100</position>
<input>
<ID>J</ID>931 </input>
<input>
<ID>K</ID>931 </input>
<output>
<ID>Q</ID>937 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>910</ID>
<type>BB_CLOCK</type>
<position>-590,-40.5</position>
<output>
<ID>CLK</ID>895 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 3</lparam></gate>
<gate>
<ID>911</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-356,-100</position>
<input>
<ID>J</ID>932 </input>
<input>
<ID>K</ID>932 </input>
<output>
<ID>Q</ID>938 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>912</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-344,-114.5</position>
<input>
<ID>IN_0</ID>933 </input>
<input>
<ID>IN_1</ID>934 </input>
<input>
<ID>IN_2</ID>936 </input>
<input>
<ID>IN_3</ID>935 </input>
<input>
<ID>IN_4</ID>937 </input>
<input>
<ID>IN_5</ID>938 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>913</ID>
<type>AA_AND2</type>
<position>-542.5,-16.5</position>
<input>
<ID>IN_0</ID>916 </input>
<input>
<ID>IN_1</ID>918 </input>
<output>
<ID>OUT</ID>912 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>914</ID>
<type>AA_AND2</type>
<position>-414,-89.5</position>
<input>
<ID>IN_0</ID>933 </input>
<input>
<ID>IN_1</ID>934 </input>
<output>
<ID>OUT</ID>929 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>915</ID>
<type>AA_AND2</type>
<position>-397,-90.5</position>
<input>
<ID>IN_0</ID>929 </input>
<input>
<ID>IN_1</ID>936 </input>
<output>
<ID>OUT</ID>930 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>916</ID>
<type>AA_AND2</type>
<position>-525.5,-17.5</position>
<input>
<ID>IN_0</ID>912 </input>
<input>
<ID>IN_1</ID>920 </input>
<output>
<ID>OUT</ID>913 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>917</ID>
<type>AA_AND2</type>
<position>-382,-91.5</position>
<input>
<ID>IN_0</ID>930 </input>
<input>
<ID>IN_1</ID>935 </input>
<output>
<ID>OUT</ID>931 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>918</ID>
<type>AA_AND2</type>
<position>-364.5,-92.5</position>
<input>
<ID>IN_0</ID>931 </input>
<input>
<ID>IN_1</ID>937 </input>
<output>
<ID>OUT</ID>932 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>919</ID>
<type>AA_AND2</type>
<position>-510.5,-18.5</position>
<input>
<ID>IN_0</ID>913 </input>
<input>
<ID>IN_1</ID>919 </input>
<output>
<ID>OUT</ID>914 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>920</ID>
<type>BA_NAND4</type>
<position>-342.5,-89.5</position>
<input>
<ID>IN_0</ID>936 </input>
<input>
<ID>IN_1</ID>935 </input>
<input>
<ID>IN_2</ID>937 </input>
<input>
<ID>IN_3</ID>938 </input>
<output>
<ID>OUT</ID>905 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>921</ID>
<type>AE_DFF_LOW</type>
<position>-425.5,-135</position>
<input>
<ID>IN_0</ID>933 </input>
<output>
<ID>OUT_0</ID>939 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>922</ID>
<type>AA_AND2</type>
<position>-493,-19.5</position>
<input>
<ID>IN_0</ID>914 </input>
<input>
<ID>IN_1</ID>921 </input>
<output>
<ID>OUT</ID>915 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>923</ID>
<type>AE_DFF_LOW</type>
<position>-409,-135</position>
<input>
<ID>IN_0</ID>934 </input>
<output>
<ID>OUT_0</ID>940 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>924</ID>
<type>AE_DFF_LOW</type>
<position>-394.5,-135</position>
<input>
<ID>IN_0</ID>936 </input>
<output>
<ID>OUT_0</ID>941 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>925</ID>
<type>BA_NAND4</type>
<position>-471,-16.5</position>
<input>
<ID>IN_0</ID>920 </input>
<input>
<ID>IN_1</ID>919 </input>
<input>
<ID>IN_2</ID>921 </input>
<input>
<ID>IN_3</ID>922 </input>
<output>
<ID>OUT</ID>904 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>926</ID>
<type>AE_DFF_LOW</type>
<position>-377.5,-135</position>
<input>
<ID>IN_0</ID>935 </input>
<output>
<ID>OUT_0</ID>942 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>927</ID>
<type>AE_DFF_LOW</type>
<position>-361.5,-135</position>
<input>
<ID>IN_0</ID>937 </input>
<output>
<ID>OUT_0</ID>943 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>928</ID>
<type>AE_DFF_LOW</type>
<position>-343.5,-135</position>
<input>
<ID>IN_0</ID>938 </input>
<output>
<ID>OUT_0</ID>944 </output>
<input>
<ID>clear</ID>899 </input>
<input>
<ID>clock</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>929</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-323.5,-144.5</position>
<input>
<ID>IN_0</ID>939 </input>
<input>
<ID>IN_1</ID>940 </input>
<input>
<ID>IN_2</ID>941 </input>
<input>
<ID>IN_3</ID>942 </input>
<input>
<ID>IN_4</ID>943 </input>
<input>
<ID>IN_5</ID>944 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>930</ID>
<type>AA_INVERTER</type>
<position>-436,-42</position>
<input>
<ID>IN_0</ID>903 </input>
<output>
<ID>OUT_0</ID>946 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>931</ID>
<type>AE_DFF_LOW</type>
<position>-554,-62</position>
<input>
<ID>IN_0</ID>916 </input>
<output>
<ID>OUT_0</ID>923 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>932</ID>
<type>AE_DFF_LOW</type>
<position>-537.5,-62</position>
<input>
<ID>IN_0</ID>918 </input>
<output>
<ID>OUT_0</ID>924 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>933</ID>
<type>AE_DFF_LOW</type>
<position>-523,-62</position>
<input>
<ID>IN_0</ID>920 </input>
<output>
<ID>OUT_0</ID>925 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>934</ID>
<type>AE_DFF_LOW</type>
<position>-506,-62</position>
<input>
<ID>IN_0</ID>919 </input>
<output>
<ID>OUT_0</ID>926 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>935</ID>
<type>AE_DFF_LOW</type>
<position>-490,-62</position>
<input>
<ID>IN_0</ID>921 </input>
<output>
<ID>OUT_0</ID>927 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>936</ID>
<type>AE_DFF_LOW</type>
<position>-472,-62</position>
<input>
<ID>IN_0</ID>922 </input>
<output>
<ID>OUT_0</ID>928 </output>
<input>
<ID>clear</ID>903 </input>
<input>
<ID>clock</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>937</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-452,-71.5</position>
<input>
<ID>IN_0</ID>923 </input>
<input>
<ID>IN_1</ID>924 </input>
<input>
<ID>IN_2</ID>925 </input>
<input>
<ID>IN_3</ID>926 </input>
<input>
<ID>IN_4</ID>927 </input>
<input>
<ID>IN_5</ID>928 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>938</ID>
<type>AA_AND2</type>
<position>-589.5,-31</position>
<input>
<ID>IN_0</ID>826 </input>
<input>
<ID>IN_1</ID>833 </input>
<output>
<ID>OUT</ID>945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>939</ID>
<type>AE_DFF_LOW</type>
<position>-645.5,-198</position>
<input>
<ID>IN_0</ID>828 </input>
<output>
<ID>OUTINV_0</ID>834 </output>
<output>
<ID>OUT_0</ID>832 </output>
<input>
<ID>clock</ID>830 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>940</ID>
<type>AI_XOR2</type>
<position>-101,-418</position>
<input>
<ID>IN_0</ID>939 </input>
<input>
<ID>IN_1</ID>842 </input>
<output>
<ID>OUT</ID>805 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>941</ID>
<type>AA_TOGGLE</type>
<position>-658,-196</position>
<output>
<ID>OUT_0</ID>828 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>942</ID>
<type>AI_XOR2</type>
<position>-87.5,-418</position>
<input>
<ID>IN_0</ID>940 </input>
<input>
<ID>IN_1</ID>860 </input>
<output>
<ID>OUT</ID>806 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>943</ID>
<type>AI_XOR2</type>
<position>-74.5,-418</position>
<input>
<ID>IN_0</ID>941 </input>
<input>
<ID>IN_1</ID>861 </input>
<output>
<ID>OUT</ID>807 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>944</ID>
<type>AA_AND2</type>
<position>-629,-187</position>
<input>
<ID>IN_0</ID>832 </input>
<input>
<ID>IN_1</ID>831 </input>
<output>
<ID>OUT</ID>833 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>945</ID>
<type>AI_XOR2</type>
<position>-61.5,-418</position>
<input>
<ID>IN_0</ID>942 </input>
<input>
<ID>IN_1</ID>862 </input>
<output>
<ID>OUT</ID>808 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>946</ID>
<type>AA_LABEL</type>
<position>-662,-186.5</position>
<gparam>LABEL_TEXT On/Off Switch</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>947</ID>
<type>AI_XOR2</type>
<position>-49,-418.5</position>
<input>
<ID>IN_0</ID>943 </input>
<input>
<ID>IN_1</ID>863 </input>
<output>
<ID>OUT</ID>809 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>948</ID>
<type>AI_XOR2</type>
<position>-36.5,-418.5</position>
<input>
<ID>IN_0</ID>944 </input>
<input>
<ID>IN_1</ID>864 </input>
<output>
<ID>OUT</ID>810 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>949</ID>
<type>AE_SMALL_INVERTER</type>
<position>-635,-199</position>
<input>
<ID>IN_0</ID>834 </input>
<output>
<ID>OUT_0</ID>835 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>805</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-101,-424.5,-101,-421</points>
<connection>
<GID>940</GID>
<name>OUT</name></connection>
<intersection>-424.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-101,-424.5,-100,-424.5</points>
<connection>
<GID>788</GID>
<name>IN_0</name></connection>
<intersection>-101 0</intersection></hsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,-425,-87.5,-421</points>
<connection>
<GID>942</GID>
<name>OUT</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-425,-84,-425</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>-87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,-425,-74.5,-421</points>
<connection>
<GID>943</GID>
<name>OUT</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74.5,-425,-70.5,-425</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>-74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-425,-58.5,-421</points>
<intersection>-425 1</intersection>
<intersection>-421 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,-425,-55.5,-425</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-61.5,-421,-58.5,-421</points>
<connection>
<GID>945</GID>
<name>OUT</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-423.5,-49,-421.5</points>
<connection>
<GID>947</GID>
<name>OUT</name></connection>
<intersection>-423.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-423.5,-45,-423.5</points>
<intersection>-49 0</intersection>
<intersection>-45 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-45,-425,-45,-423.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>-423.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-423.5,-36.5,-421.5</points>
<connection>
<GID>948</GID>
<name>OUT</name></connection>
<intersection>-423.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-423.5,-32,-423.5</points>
<intersection>-36.5 0</intersection>
<intersection>-32 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-32,-425,-32,-423.5</points>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>-423.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90,-432.5,-90,-424.5</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>-424.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94,-424.5,-90,-424.5</points>
<connection>
<GID>788</GID>
<name>OUT_0</name></connection>
<intersection>-90 0</intersection></hsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,-432.5,-75,-425</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,-425,-75,-425</points>
<connection>
<GID>789</GID>
<name>OUT_0</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-432.5,-60,-425</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-425,-60,-425</points>
<connection>
<GID>790</GID>
<name>OUT_0</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,-432,-48.5,-425</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-425,-48.5,-425</points>
<connection>
<GID>791</GID>
<name>OUT_0</name></connection>
<intersection>-48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-432.5,-35.5,-425</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-425,-35.5,-425</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>816</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-432,-22.5,-425</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-425,-22.5,-425</points>
<connection>
<GID>793</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>817</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90,-442,-90,-436.5</points>
<connection>
<GID>794</GID>
<name>OUT_0</name></connection>
<intersection>-442 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-75,-448,-75,-442</points>
<connection>
<GID>800</GID>
<name>IN_3</name></connection>
<intersection>-442 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-90,-442,-75,-442</points>
<intersection>-90 0</intersection>
<intersection>-75 1</intersection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,-441.5,-75,-436.5</points>
<connection>
<GID>795</GID>
<name>OUT_0</name></connection>
<intersection>-441.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-73,-448,-73,-441.5</points>
<connection>
<GID>800</GID>
<name>IN_2</name></connection>
<intersection>-441.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-75,-441.5,-73,-441.5</points>
<intersection>-75 0</intersection>
<intersection>-73 1</intersection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-442,-60,-436.5</points>
<connection>
<GID>796</GID>
<name>OUT_0</name></connection>
<intersection>-442 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-71,-448,-71,-442</points>
<connection>
<GID>800</GID>
<name>IN_1</name></connection>
<intersection>-442 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-71,-442,-60,-442</points>
<intersection>-71 1</intersection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,-443,-48.5,-436</points>
<connection>
<GID>797</GID>
<name>OUT_0</name></connection>
<intersection>-443 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-69,-448,-69,-443</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<intersection>-443 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-69,-443,-48.5,-443</points>
<intersection>-69 1</intersection>
<intersection>-48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-441.5,-35.5,-436.5</points>
<connection>
<GID>798</GID>
<name>OUT_0</name></connection>
<intersection>-441.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-36.5,-447,-36.5,-441.5</points>
<connection>
<GID>801</GID>
<name>IN_1</name></connection>
<intersection>-441.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,-441.5,-35.5,-441.5</points>
<intersection>-36.5 1</intersection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-441.5,-22.5,-436</points>
<connection>
<GID>799</GID>
<name>OUT_0</name></connection>
<intersection>-441.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-34.5,-447,-34.5,-441.5</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<intersection>-441.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-441.5,-22.5,-441.5</points>
<intersection>-34.5 1</intersection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>823</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,-457,-72,-454</points>
<connection>
<GID>800</GID>
<name>OUT</name></connection>
<intersection>-457 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-57.5,-460,-57.5,-457</points>
<connection>
<GID>802</GID>
<name>IN_1</name></connection>
<intersection>-457 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-72,-457,-57.5,-457</points>
<intersection>-72 0</intersection>
<intersection>-57.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-456.5,-35.5,-453</points>
<connection>
<GID>801</GID>
<name>OUT</name></connection>
<intersection>-456.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-55.5,-460,-55.5,-456.5</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<intersection>-456.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-456.5,-35.5,-456.5</points>
<intersection>-55.5 1</intersection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-582,-11.5,-582,-7</points>
<connection>
<GID>803</GID>
<name>IN_1</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-591.5,-7,-582,-7</points>
<connection>
<GID>899</GID>
<name>OUT_0</name></connection>
<intersection>-582 0</intersection></hsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-593.5,-30,-593.5,-17.5</points>
<intersection>-30 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-593.5,-30,-592.5,-30</points>
<connection>
<GID>938</GID>
<name>IN_0</name></connection>
<intersection>-593.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-593.5,-17.5,-581,-17.5</points>
<connection>
<GID>803</GID>
<name>OUT</name></connection>
<intersection>-593.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-466,-4,-2.5</points>
<intersection>-466 4</intersection>
<intersection>-2.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-580,-2.5,-4,-2.5</points>
<intersection>-580 5</intersection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-56.5,-466,-4,-466</points>
<connection>
<GID>802</GID>
<name>OUT</name></connection>
<intersection>-4 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-580,-11.5,-580,-2.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>-2.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-656,-196,-648.5,-196</points>
<connection>
<GID>939</GID>
<name>IN_0</name></connection>
<connection>
<GID>941</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-606.5,-198,-598.5,-198</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<connection>
<GID>808</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-602.5,-206.5,-602.5,-201</points>
<intersection>-206.5 2</intersection>
<intersection>-201 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-602.5,-201,-598.5,-201</points>
<connection>
<GID>805</GID>
<name>clock</name></connection>
<intersection>-602.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-648.5,-206.5,-602.5,-206.5</points>
<intersection>-648.5 3</intersection>
<intersection>-606.5 4</intersection>
<intersection>-602.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-648.5,-206.5,-648.5,-199</points>
<connection>
<GID>939</GID>
<name>clock</name></connection>
<intersection>-206.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-606.5,-206.5,-606.5,-203.5</points>
<connection>
<GID>806</GID>
<name>CLK</name></connection>
<intersection>-206.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-628,-210,-628,-190</points>
<connection>
<GID>944</GID>
<name>IN_1</name></connection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-628,-210,-592.5,-210</points>
<intersection>-628 0</intersection>
<intersection>-592.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-592.5,-210,-592.5,-201</points>
<connection>
<GID>805</GID>
<name>OUTINV_0</name></connection>
<intersection>-210 1</intersection></vsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-630,-196,-630,-190</points>
<connection>
<GID>944</GID>
<name>IN_0</name></connection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-642.5,-196,-630,-196</points>
<connection>
<GID>939</GID>
<name>OUT_0</name></connection>
<intersection>-630 0</intersection></hsegment></shape></wire>
<wire>
<ID>833</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-629,-184,-629,-32</points>
<connection>
<GID>944</GID>
<name>OUT</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-629,-32,-592.5,-32</points>
<connection>
<GID>938</GID>
<name>IN_1</name></connection>
<intersection>-629 0</intersection></hsegment></shape></wire>
<wire>
<ID>834</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-642.5,-199,-637,-199</points>
<connection>
<GID>939</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>949</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-595.5,-239,-595.5,-204</points>
<connection>
<GID>805</GID>
<name>clear</name></connection>
<intersection>-239 3</intersection>
<intersection>-211.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-633,-211.5,-595.5,-211.5</points>
<intersection>-633 2</intersection>
<intersection>-595.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-633,-211.5,-633,-199</points>
<connection>
<GID>949</GID>
<name>OUT_0</name></connection>
<intersection>-211.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-595.5,-239,-580,-239</points>
<connection>
<GID>839</GID>
<name>clear</name></connection>
<intersection>-595.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>836</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-291.5,-256.5,-291.5,-201</points>
<intersection>-256.5 2</intersection>
<intersection>-201 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-296.5,-201,-291.5,-201</points>
<connection>
<GID>810</GID>
<name>OUT</name></connection>
<intersection>-291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-516.5,-256.5,-291.5,-256.5</points>
<intersection>-516.5 15</intersection>
<intersection>-467 14</intersection>
<intersection>-441 10</intersection>
<intersection>-411 18</intersection>
<intersection>-372.5 16</intersection>
<intersection>-324 17</intersection>
<intersection>-291.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-441,-256.5,-441,-230.5</points>
<connection>
<GID>815</GID>
<name>clear</name></connection>
<intersection>-256.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-467,-256.5,-467,-231</points>
<connection>
<GID>813</GID>
<name>clear</name></connection>
<intersection>-256.5 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-516.5,-256.5,-516.5,-230.5</points>
<connection>
<GID>812</GID>
<name>clear</name></connection>
<intersection>-256.5 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-372.5,-256.5,-372.5,-233</points>
<connection>
<GID>817</GID>
<name>clear</name></connection>
<intersection>-256.5 2</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-324,-256.5,-324,-233.5</points>
<connection>
<GID>818</GID>
<name>clear</name></connection>
<intersection>-256.5 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-411,-256.5,-411,-231</points>
<connection>
<GID>816</GID>
<name>clear</name></connection>
<intersection>-256.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-507.5,-269,-507.5,-218.5</points>
<intersection>-269 8</intersection>
<intersection>-263 5</intersection>
<intersection>-253.5 3</intersection>
<intersection>-224.5 2</intersection>
<intersection>-218.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-507.5,-218.5,-503,-218.5</points>
<connection>
<GID>820</GID>
<name>IN_1</name></connection>
<intersection>-507.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-513.5,-224.5,-507.5,-224.5</points>
<connection>
<GID>812</GID>
<name>Q</name></connection>
<intersection>-507.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-507.5,-253.5,-304.5,-253.5</points>
<connection>
<GID>838</GID>
<name>IN_0</name></connection>
<intersection>-507.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-507.5,-263,-488.5,-263</points>
<intersection>-507.5 0</intersection>
<intersection>-488.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-488.5,-295.5,-488.5,-263</points>
<connection>
<GID>859</GID>
<name>IN_0</name></connection>
<intersection>-263 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-507.5,-269,-501.5,-269</points>
<connection>
<GID>811</GID>
<name>IN_0</name></connection>
<intersection>-507.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-511.5,-234,-511.5,-228.5</points>
<intersection>-234 3</intersection>
<intersection>-228.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-513.5,-228.5,-511.5,-228.5</points>
<connection>
<GID>812</GID>
<name>nQ</name></connection>
<intersection>-511.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-511.5,-234,-504,-234</points>
<connection>
<GID>821</GID>
<name>IN_0</name></connection>
<intersection>-511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-493,-226,-493,-216.5</points>
<intersection>-226 1</intersection>
<intersection>-217.5 2</intersection>
<intersection>-216.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-493,-226,-489,-226</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>-493 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-497,-217.5,-493,-217.5</points>
<connection>
<GID>820</GID>
<name>OUT</name></connection>
<intersection>-493 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-493,-216.5,-462,-216.5</points>
<connection>
<GID>822</GID>
<name>IN_0</name></connection>
<intersection>-493 0</intersection></hsegment></shape></wire>
<wire>
<ID>840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-492.5,-237,-492.5,-228</points>
<intersection>-237 2</intersection>
<intersection>-235 3</intersection>
<intersection>-228 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-492.5,-228,-489,-228</points>
<connection>
<GID>831</GID>
<name>IN_1</name></connection>
<intersection>-492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-492.5,-237,-459.5,-237</points>
<connection>
<GID>823</GID>
<name>IN_1</name></connection>
<intersection>-492.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-498,-235,-492.5,-235</points>
<connection>
<GID>821</GID>
<name>OUT</name></connection>
<intersection>-492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-463,-295,-463,-218.5</points>
<intersection>-295 9</intersection>
<intersection>-268.5 5</intersection>
<intersection>-252.5 3</intersection>
<intersection>-225 2</intersection>
<intersection>-218.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-463,-218.5,-462,-218.5</points>
<connection>
<GID>822</GID>
<name>IN_1</name></connection>
<intersection>-463 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-464,-225,-463,-225</points>
<connection>
<GID>813</GID>
<name>Q</name></connection>
<intersection>-463 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-463,-252.5,-304.5,-252.5</points>
<connection>
<GID>838</GID>
<name>IN_1</name></connection>
<intersection>-463 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-463,-268.5,-458.5,-268.5</points>
<connection>
<GID>814</GID>
<name>IN_0</name></connection>
<intersection>-463 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-476,-295,-463,-295</points>
<intersection>-476 10</intersection>
<intersection>-463 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-476,-296.5,-476,-295</points>
<connection>
<GID>860</GID>
<name>IN_0</name></connection>
<intersection>-295 9</intersection></vsegment></shape></wire>
<wire>
<ID>842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-492.5,-379,-492.5,-269</points>
<intersection>-379 2</intersection>
<intersection>-284 5</intersection>
<intersection>-269 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-495.5,-269,-492.5,-269</points>
<connection>
<GID>811</GID>
<name>OUT_0</name></connection>
<intersection>-492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-492.5,-379,-102,-379</points>
<intersection>-492.5 0</intersection>
<intersection>-102 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-492.5,-284,-285,-284</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>-492.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-102,-415,-102,-379</points>
<connection>
<GID>940</GID>
<name>IN_1</name></connection>
<intersection>-379 2</intersection></vsegment></shape></wire>
<wire>
<ID>843</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-454.5,-218,-454.5,-217.5</points>
<intersection>-218 2</intersection>
<intersection>-217.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-456,-217.5,-454.5,-217.5</points>
<connection>
<GID>822</GID>
<name>OUT</name></connection>
<intersection>-454.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-454.5,-218,-432.5,-218</points>
<connection>
<GID>824</GID>
<name>IN_0</name></connection>
<intersection>-454.5 0</intersection>
<intersection>-452.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-452.5,-225,-452.5,-218</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<intersection>-218 2</intersection></vsegment></shape></wire>
<wire>
<ID>844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-461.5,-235,-461.5,-229</points>
<intersection>-235 2</intersection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-464,-229,-461.5,-229</points>
<connection>
<GID>813</GID>
<name>nQ</name></connection>
<intersection>-461.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-461.5,-235,-459.5,-235</points>
<connection>
<GID>823</GID>
<name>IN_0</name></connection>
<intersection>-461.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-453,-238.5,-453,-227</points>
<intersection>-238.5 3</intersection>
<intersection>-236 1</intersection>
<intersection>-227 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-453.5,-236,-453,-236</points>
<connection>
<GID>823</GID>
<name>OUT</name></connection>
<intersection>-453 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-453,-227,-452.5,-227</points>
<connection>
<GID>833</GID>
<name>IN_1</name></connection>
<intersection>-453 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-453,-238.5,-430,-238.5</points>
<connection>
<GID>825</GID>
<name>IN_1</name></connection>
<intersection>-453 0</intersection></hsegment></shape></wire>
<wire>
<ID>846</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-436,-295.5,-436,-198</points>
<intersection>-295.5 13</intersection>
<intersection>-268.5 9</intersection>
<intersection>-251.5 2</intersection>
<intersection>-224.5 1</intersection>
<intersection>-220 5</intersection>
<intersection>-198 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-438,-224.5,-436,-224.5</points>
<connection>
<GID>815</GID>
<name>Q</name></connection>
<intersection>-436 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-436,-251.5,-304.5,-251.5</points>
<connection>
<GID>838</GID>
<name>IN_2</name></connection>
<intersection>-436 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-436,-220,-432.5,-220</points>
<connection>
<GID>824</GID>
<name>IN_1</name></connection>
<intersection>-436 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-436,-198,-302.5,-198</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-436 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-436,-268.5,-429,-268.5</points>
<connection>
<GID>819</GID>
<name>IN_0</name></connection>
<intersection>-436 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-436,-295.5,-412,-295.5</points>
<connection>
<GID>861</GID>
<name>IN_0</name></connection>
<intersection>-436 0</intersection></hsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-426.5,-219,-406,-219</points>
<connection>
<GID>824</GID>
<name>OUT</name></connection>
<connection>
<GID>826</GID>
<name>IN_0</name></connection>
<intersection>-424 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-424,-225.5,-424,-219</points>
<connection>
<GID>834</GID>
<name>IN_0</name></connection>
<intersection>-219 1</intersection></vsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-424,-238.5,-424,-227.5</points>
<connection>
<GID>834</GID>
<name>IN_1</name></connection>
<connection>
<GID>825</GID>
<name>OUT</name></connection>
<intersection>-238.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-424,-238.5,-404.5,-238.5</points>
<connection>
<GID>827</GID>
<name>IN_1</name></connection>
<intersection>-424 0</intersection></hsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-434.5,-236.5,-434.5,-228.5</points>
<intersection>-236.5 2</intersection>
<intersection>-228.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-438,-228.5,-434.5,-228.5</points>
<connection>
<GID>815</GID>
<name>nQ</name></connection>
<intersection>-434.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-434.5,-236.5,-430,-236.5</points>
<connection>
<GID>825</GID>
<name>IN_0</name></connection>
<intersection>-434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>850</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-408,-268.5,-408,-200</points>
<connection>
<GID>816</GID>
<name>Q</name></connection>
<intersection>-268.5 10</intersection>
<intersection>-250.5 2</intersection>
<intersection>-221 6</intersection>
<intersection>-200 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-408,-250.5,-304.5,-250.5</points>
<connection>
<GID>838</GID>
<name>IN_3</name></connection>
<intersection>-408 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-408,-221,-406,-221</points>
<connection>
<GID>826</GID>
<name>IN_1</name></connection>
<intersection>-408 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-408,-200,-302.5,-200</points>
<connection>
<GID>810</GID>
<name>IN_1</name></connection>
<intersection>-408 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-408,-268.5,-400.5,-268.5</points>
<connection>
<GID>830</GID>
<name>IN_0</name></connection>
<intersection>-408 0</intersection>
<intersection>-405 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-405,-295.5,-405,-268.5</points>
<connection>
<GID>862</GID>
<name>IN_0</name></connection>
<intersection>-268.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-407,-236.5,-407,-229</points>
<intersection>-236.5 2</intersection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-408,-229,-407,-229</points>
<connection>
<GID>816</GID>
<name>nQ</name></connection>
<intersection>-407 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-407,-236.5,-404.5,-236.5</points>
<connection>
<GID>827</GID>
<name>IN_0</name></connection>
<intersection>-407 0</intersection></hsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-397,-226,-397,-218</points>
<intersection>-226 2</intersection>
<intersection>-220 1</intersection>
<intersection>-218 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-400,-220,-397,-220</points>
<connection>
<GID>826</GID>
<name>OUT</name></connection>
<intersection>-397 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-397,-226,-395,-226</points>
<connection>
<GID>835</GID>
<name>IN_0</name></connection>
<intersection>-397 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-397,-218,-359,-218</points>
<connection>
<GID>828</GID>
<name>IN_0</name></connection>
<intersection>-397 0</intersection></hsegment></shape></wire>
<wire>
<ID>853</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-396.5,-237.5,-396.5,-228</points>
<intersection>-237.5 1</intersection>
<intersection>-228 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-398.5,-237.5,-358.5,-237.5</points>
<connection>
<GID>827</GID>
<name>OUT</name></connection>
<connection>
<GID>829</GID>
<name>IN_1</name></connection>
<intersection>-396.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-396.5,-228,-395,-228</points>
<connection>
<GID>835</GID>
<name>IN_1</name></connection>
<intersection>-396.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-364.5,-295,-364.5,-202</points>
<intersection>-295 14</intersection>
<intersection>-268.5 9</intersection>
<intersection>-249.5 3</intersection>
<intersection>-227 1</intersection>
<intersection>-220 10</intersection>
<intersection>-202 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-369.5,-227,-364.5,-227</points>
<connection>
<GID>817</GID>
<name>Q</name></connection>
<intersection>-364.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-364.5,-249.5,-304.5,-249.5</points>
<connection>
<GID>838</GID>
<name>IN_4</name></connection>
<intersection>-364.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-364.5,-202,-302.5,-202</points>
<connection>
<GID>810</GID>
<name>IN_2</name></connection>
<intersection>-364.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-364.5,-268.5,-354.5,-268.5</points>
<connection>
<GID>832</GID>
<name>IN_0</name></connection>
<intersection>-364.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-364.5,-220,-359,-220</points>
<connection>
<GID>828</GID>
<name>IN_1</name></connection>
<intersection>-364.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-364.5,-295,-347.5,-295</points>
<connection>
<GID>863</GID>
<name>IN_0</name></connection>
<intersection>-364.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>855</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-367,-235.5,-367,-231</points>
<intersection>-235.5 2</intersection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-369.5,-231,-367,-231</points>
<connection>
<GID>817</GID>
<name>nQ</name></connection>
<intersection>-367 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-367,-235.5,-358.5,-235.5</points>
<connection>
<GID>829</GID>
<name>IN_0</name></connection>
<intersection>-367 0</intersection></hsegment></shape></wire>
<wire>
<ID>856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-352,-226.5,-352,-219</points>
<intersection>-226.5 2</intersection>
<intersection>-219 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-353,-219,-352,-219</points>
<connection>
<GID>828</GID>
<name>OUT</name></connection>
<intersection>-352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-352,-226.5,-351,-226.5</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>-352 0</intersection></hsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-352,-236.5,-352,-228.5</points>
<intersection>-236.5 1</intersection>
<intersection>-228.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-352.5,-236.5,-352,-236.5</points>
<connection>
<GID>829</GID>
<name>OUT</name></connection>
<intersection>-352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-352,-228.5,-351,-228.5</points>
<connection>
<GID>836</GID>
<name>IN_1</name></connection>
<intersection>-352 0</intersection></hsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-545,-246,-327,-246</points>
<intersection>-545 16</intersection>
<intersection>-527.5 13</intersection>
<intersection>-470.5 12</intersection>
<intersection>-445 6</intersection>
<intersection>-417 7</intersection>
<intersection>-379 11</intersection>
<intersection>-327 28</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-445,-246,-445,-226.5</points>
<intersection>-246 1</intersection>
<intersection>-226.5 19</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-417,-246,-417,-227</points>
<intersection>-246 1</intersection>
<intersection>-227 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-379,-246,-379,-229</points>
<intersection>-246 1</intersection>
<intersection>-229 18</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-470.5,-246,-470.5,-227</points>
<intersection>-246 1</intersection>
<intersection>-227 22</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-527.5,-246,-527.5,-226.5</points>
<intersection>-246 1</intersection>
<intersection>-226.5 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-417,-227,-414,-227</points>
<connection>
<GID>816</GID>
<name>clock</name></connection>
<intersection>-417 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-527.5,-226.5,-519.5,-226.5</points>
<connection>
<GID>812</GID>
<name>clock</name></connection>
<intersection>-527.5 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-545,-275.5,-545,-246</points>
<intersection>-275.5 17</intersection>
<intersection>-246.5 37</intersection>
<intersection>-246 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-545,-275.5,-306.5,-275.5</points>
<intersection>-545 16</intersection>
<intersection>-501.5 34</intersection>
<intersection>-458.5 25</intersection>
<intersection>-429 26</intersection>
<intersection>-400.5 24</intersection>
<intersection>-355.5 23</intersection>
<intersection>-306.5 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-379,-229,-375.5,-229</points>
<connection>
<GID>817</GID>
<name>clock</name></connection>
<intersection>-379 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-445,-226.5,-444,-226.5</points>
<connection>
<GID>815</GID>
<name>clock</name></connection>
<intersection>-445 6</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-470.5,-227,-470,-227</points>
<connection>
<GID>813</GID>
<name>clock</name></connection>
<intersection>-470.5 12</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-355.5,-275.5,-355.5,-271.5</points>
<intersection>-275.5 17</intersection>
<intersection>-271.5 36</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-400.5,-275.5,-400.5,-271.5</points>
<connection>
<GID>830</GID>
<name>clock</name></connection>
<intersection>-275.5 17</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>-458.5,-275.5,-458.5,-271.5</points>
<connection>
<GID>814</GID>
<name>clock</name></connection>
<intersection>-275.5 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-429,-275.5,-429,-271.5</points>
<connection>
<GID>819</GID>
<name>clock</name></connection>
<intersection>-275.5 17</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-327,-246,-327,-229.5</points>
<connection>
<GID>818</GID>
<name>clock</name></connection>
<intersection>-246 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-501.5,-275.5,-501.5,-272</points>
<connection>
<GID>811</GID>
<name>clock</name></connection>
<intersection>-275.5 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>-306.5,-275.5,-306.5,-272</points>
<connection>
<GID>837</GID>
<name>clock</name></connection>
<intersection>-275.5 17</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>-355.5,-271.5,-354.5,-271.5</points>
<connection>
<GID>832</GID>
<name>clock</name></connection>
<intersection>-355.5 23</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-586,-246.5,-545,-246.5</points>
<connection>
<GID>844</GID>
<name>OUT</name></connection>
<intersection>-583.5 38</intersection>
<intersection>-545 16</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>-583.5,-246.5,-583.5,-236</points>
<intersection>-246.5 37</intersection>
<intersection>-236 39</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-583.5,-236,-583,-236</points>
<connection>
<GID>839</GID>
<name>clock</name></connection>
<intersection>-583.5 38</intersection></hsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-312,-294.5,-312,-204</points>
<intersection>-294.5 9</intersection>
<intersection>-269 13</intersection>
<intersection>-248.5 2</intersection>
<intersection>-227.5 11</intersection>
<intersection>-204 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-312,-248.5,-304.5,-248.5</points>
<connection>
<GID>838</GID>
<name>IN_5</name></connection>
<intersection>-312 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-312,-204,-302.5,-204</points>
<connection>
<GID>810</GID>
<name>IN_3</name></connection>
<intersection>-312 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-342,-294.5,-312,-294.5</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<intersection>-312 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-321,-227.5,-312,-227.5</points>
<connection>
<GID>818</GID>
<name>Q</name></connection>
<intersection>-312 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-312,-269,-306.5,-269</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<intersection>-312 0</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-451,-370.5,-451,-268.5</points>
<intersection>-370.5 7</intersection>
<intersection>-268.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-452.5,-268.5,-451,-268.5</points>
<connection>
<GID>814</GID>
<name>OUT_0</name></connection>
<intersection>-451 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-451,-370.5,-88.5,-370.5</points>
<intersection>-451 3</intersection>
<intersection>-285 10</intersection>
<intersection>-88.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88.5,-415,-88.5,-370.5</points>
<connection>
<GID>942</GID>
<name>IN_1</name></connection>
<intersection>-370.5 7</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-285,-370.5,-285,-283</points>
<connection>
<GID>841</GID>
<name>IN_1</name></connection>
<intersection>-370.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-421.5,-357.5,-75.5,-357.5</points>
<intersection>-421.5 3</intersection>
<intersection>-75.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-421.5,-357.5,-421.5,-268.5</points>
<intersection>-357.5 1</intersection>
<intersection>-282 7</intersection>
<intersection>-268.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-423,-268.5,-421.5,-268.5</points>
<connection>
<GID>819</GID>
<name>OUT_0</name></connection>
<intersection>-421.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-421.5,-282,-285,-282</points>
<connection>
<GID>841</GID>
<name>IN_2</name></connection>
<intersection>-421.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-75.5,-415,-75.5,-357.5</points>
<connection>
<GID>943</GID>
<name>IN_1</name></connection>
<intersection>-357.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-394.5,-350.5,-62.5,-350.5</points>
<intersection>-394.5 3</intersection>
<intersection>-62.5 12</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-394.5,-350.5,-394.5,-268.5</points>
<connection>
<GID>830</GID>
<name>OUT_0</name></connection>
<intersection>-350.5 1</intersection>
<intersection>-281 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-394.5,-281,-285,-281</points>
<connection>
<GID>841</GID>
<name>IN_3</name></connection>
<intersection>-394.5 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-62.5,-415,-62.5,-350.5</points>
<connection>
<GID>945</GID>
<name>IN_1</name></connection>
<intersection>-350.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>863</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-336.5,-343,-336.5,-268.5</points>
<intersection>-343 2</intersection>
<intersection>-280 5</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-348.5,-268.5,-336.5,-268.5</points>
<connection>
<GID>832</GID>
<name>OUT_0</name></connection>
<intersection>-336.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-336.5,-343,-50,-343</points>
<intersection>-336.5 0</intersection>
<intersection>-50 7</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-336.5,-280,-285,-280</points>
<connection>
<GID>841</GID>
<name>IN_4</name></connection>
<intersection>-336.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-50,-415.5,-50,-343</points>
<connection>
<GID>947</GID>
<name>IN_1</name></connection>
<intersection>-343 2</intersection></vsegment></shape></wire>
<wire>
<ID>864</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-293.5,-337,-293.5,-269</points>
<intersection>-337 7</intersection>
<intersection>-279 10</intersection>
<intersection>-269 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-300.5,-269,-293.5,-269</points>
<connection>
<GID>837</GID>
<name>OUT_0</name></connection>
<intersection>-293.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-293.5,-337,-37.5,-337</points>
<intersection>-293.5 3</intersection>
<intersection>-37.5 12</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-293.5,-279,-285,-279</points>
<connection>
<GID>841</GID>
<name>IN_5</name></connection>
<intersection>-293.5 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-37.5,-415.5,-37.5,-337</points>
<connection>
<GID>948</GID>
<name>IN_1</name></connection>
<intersection>-337 7</intersection></vsegment></shape></wire>
<wire>
<ID>865</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-522.5,-224.5,-522.5,-212</points>
<intersection>-224.5 8</intersection>
<intersection>-212 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-531,-212,-522.5,-212</points>
<intersection>-531 9</intersection>
<intersection>-522.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-522.5,-224.5,-519.5,-224.5</points>
<connection>
<GID>812</GID>
<name>J</name></connection>
<intersection>-522.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-531,-212.5,-531,-200.5</points>
<connection>
<GID>852</GID>
<name>IN_0</name></connection>
<intersection>-212 6</intersection>
<intersection>-200.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-572,-200.5,-531,-200.5</points>
<intersection>-572 14</intersection>
<intersection>-531 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-572,-204,-572,-200.5</points>
<intersection>-204 15</intersection>
<intersection>-200.5 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-582.5,-204,-572,-204</points>
<connection>
<GID>867</GID>
<name>OUT</name></connection>
<intersection>-572 14</intersection></hsegment></shape></wire>
<wire>
<ID>866</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-537.5,-205,-339.5,-205</points>
<intersection>-537.5 7</intersection>
<intersection>-482 6</intersection>
<intersection>-445.5 10</intersection>
<intersection>-417 12</intersection>
<intersection>-387 14</intersection>
<intersection>-339.5 16</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-482,-210,-482,-205</points>
<connection>
<GID>853</GID>
<name>IN_1</name></connection>
<intersection>-205 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-537.5,-212,-537.5,-205</points>
<intersection>-212 20</intersection>
<intersection>-205 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-445.5,-209.5,-445.5,-205</points>
<connection>
<GID>854</GID>
<name>IN_1</name></connection>
<intersection>-205 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-417,-210,-417,-205</points>
<connection>
<GID>855</GID>
<name>IN_1</name></connection>
<intersection>-205 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-387,-210,-387,-205</points>
<connection>
<GID>856</GID>
<name>IN_1</name></connection>
<intersection>-205 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-339.5,-208,-339.5,-205</points>
<connection>
<GID>857</GID>
<name>IN_1</name></connection>
<intersection>-205 4</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-568,-212,-533,-212</points>
<intersection>-568 23</intersection>
<intersection>-537.5 7</intersection>
<intersection>-533 26</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-568,-347.5,-568,-212</points>
<intersection>-347.5 24</intersection>
<intersection>-212 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-568,-347.5,-504,-347.5</points>
<intersection>-568 23</intersection>
<intersection>-504 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-504,-347.5,-504,-346.5</points>
<connection>
<GID>858</GID>
<name>OUT</name></connection>
<intersection>-347.5 24</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-533,-212.5,-533,-212</points>
<connection>
<GID>852</GID>
<name>IN_1</name></connection>
<intersection>-212 20</intersection></vsegment></shape></wire>
<wire>
<ID>867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-532,-228.5,-532,-218.5</points>
<connection>
<GID>852</GID>
<name>OUT</name></connection>
<intersection>-228.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-532,-228.5,-519.5,-228.5</points>
<connection>
<GID>812</GID>
<name>K</name></connection>
<intersection>-532 0</intersection></hsegment></shape></wire>
<wire>
<ID>868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-483.5,-318.5,-483.5,-307</points>
<connection>
<GID>846</GID>
<name>IN_1</name></connection>
<intersection>-307 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-488.5,-307,-488.5,-301.5</points>
<connection>
<GID>859</GID>
<name>OUT_0</name></connection>
<intersection>-307 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-488.5,-307,-483.5,-307</points>
<intersection>-488.5 1</intersection>
<intersection>-483.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>869</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-481.5,-318.5,-481.5,-307</points>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>-307 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-476,-307,-476,-302.5</points>
<connection>
<GID>860</GID>
<name>OUT_0</name></connection>
<intersection>-307 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-481.5,-307,-476,-307</points>
<intersection>-481.5 0</intersection>
<intersection>-476 1</intersection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-505,-340.5,-505,-328</points>
<connection>
<GID>858</GID>
<name>IN_2</name></connection>
<intersection>-328 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-482.5,-328,-482.5,-324.5</points>
<connection>
<GID>846</GID>
<name>OUT</name></connection>
<intersection>-328 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-505,-328,-482.5,-328</points>
<intersection>-505 0</intersection>
<intersection>-482.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-407.5,-305,-407.5,-303</points>
<connection>
<GID>849</GID>
<name>IN_0</name></connection>
<intersection>-303 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-405,-303,-405,-301.5</points>
<connection>
<GID>862</GID>
<name>OUT_0</name></connection>
<intersection>-303 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-407.5,-303,-405,-303</points>
<intersection>-407.5 0</intersection>
<intersection>-405 1</intersection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-409.5,-305,-409.5,-303</points>
<connection>
<GID>849</GID>
<name>IN_1</name></connection>
<intersection>-303 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-412,-303,-412,-301.5</points>
<connection>
<GID>861</GID>
<name>OUT_0</name></connection>
<intersection>-303 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-412,-303,-409.5,-303</points>
<intersection>-412 1</intersection>
<intersection>-409.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-503,-340.5,-503,-330</points>
<connection>
<GID>858</GID>
<name>IN_1</name></connection>
<intersection>-330 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-408.5,-330,-408.5,-311</points>
<connection>
<GID>849</GID>
<name>OUT</name></connection>
<intersection>-330 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-503,-330,-408.5,-330</points>
<intersection>-503 0</intersection>
<intersection>-408.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-344.5,-303.5,-344.5,-302</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<intersection>-302 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-342,-302,-342,-300.5</points>
<connection>
<GID>864</GID>
<name>OUT_0</name></connection>
<intersection>-302 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-344.5,-302,-342,-302</points>
<intersection>-344.5 0</intersection>
<intersection>-342 1</intersection></hsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-346.5,-303.5,-346.5,-302</points>
<connection>
<GID>851</GID>
<name>IN_1</name></connection>
<intersection>-302 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-347.5,-302,-347.5,-301</points>
<connection>
<GID>863</GID>
<name>OUT_0</name></connection>
<intersection>-302 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-347.5,-302,-346.5,-302</points>
<intersection>-347.5 1</intersection>
<intersection>-346.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-501,-340.5,-501,-332.5</points>
<connection>
<GID>858</GID>
<name>IN_0</name></connection>
<intersection>-332.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-345.5,-332.5,-345.5,-309.5</points>
<connection>
<GID>851</GID>
<name>OUT</name></connection>
<intersection>-332.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-501,-332.5,-345.5,-332.5</points>
<intersection>-501 0</intersection>
<intersection>-345.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-472.5,-227,-472.5,-209.5</points>
<intersection>-227 2</intersection>
<intersection>-225 1</intersection>
<intersection>-209.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-472.5,-225,-470,-225</points>
<connection>
<GID>813</GID>
<name>J</name></connection>
<intersection>-472.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-483,-227,-472.5,-227</points>
<connection>
<GID>831</GID>
<name>OUT</name></connection>
<intersection>-472.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-480,-209.5,-472.5,-209.5</points>
<intersection>-480 4</intersection>
<intersection>-472.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-480,-210,-480,-209.5</points>
<connection>
<GID>853</GID>
<name>IN_0</name></connection>
<intersection>-209.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>878</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-481,-229,-481,-216</points>
<connection>
<GID>853</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-481,-229,-470,-229</points>
<connection>
<GID>813</GID>
<name>K</name></connection>
<intersection>-481 0</intersection></hsegment></shape></wire>
<wire>
<ID>879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-444.5,-224.5,-444.5,-215.5</points>
<connection>
<GID>854</GID>
<name>OUT</name></connection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-444.5,-224.5,-444,-224.5</points>
<connection>
<GID>815</GID>
<name>J</name></connection>
<intersection>-444.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>880</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-437,-217,-437,-209.5</points>
<intersection>-217 1</intersection>
<intersection>-209.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-446.5,-217,-437,-217</points>
<intersection>-446.5 4</intersection>
<intersection>-437 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-443.5,-209.5,-437,-209.5</points>
<connection>
<GID>854</GID>
<name>IN_0</name></connection>
<intersection>-437 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-446.5,-228.5,-446.5,-217</points>
<connection>
<GID>833</GID>
<name>OUT</name></connection>
<intersection>-228.5 6</intersection>
<intersection>-217 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-446.5,-228.5,-444,-228.5</points>
<connection>
<GID>815</GID>
<name>K</name></connection>
<intersection>-446.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>881</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-418,-217.5,-411.5,-217.5</points>
<intersection>-418 3</intersection>
<intersection>-411.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-418,-226.5,-418,-217.5</points>
<connection>
<GID>834</GID>
<name>OUT</name></connection>
<intersection>-225 7</intersection>
<intersection>-217.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-411.5,-217.5,-411.5,-210</points>
<intersection>-217.5 1</intersection>
<intersection>-210 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-415,-210,-411.5,-210</points>
<connection>
<GID>855</GID>
<name>IN_0</name></connection>
<intersection>-411.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-418,-225,-414,-225</points>
<connection>
<GID>816</GID>
<name>J</name></connection>
<intersection>-418 3</intersection></hsegment></shape></wire>
<wire>
<ID>882</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416,-229,-416,-216</points>
<connection>
<GID>855</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416,-229,-414,-229</points>
<connection>
<GID>816</GID>
<name>K</name></connection>
<intersection>-416 0</intersection></hsegment></shape></wire>
<wire>
<ID>883</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-389,-227,-375.5,-227</points>
<connection>
<GID>817</GID>
<name>J</name></connection>
<connection>
<GID>835</GID>
<name>OUT</name></connection>
<intersection>-389 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-389,-227,-389,-209</points>
<intersection>-227 1</intersection>
<intersection>-209 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-389,-209,-385,-209</points>
<intersection>-389 4</intersection>
<intersection>-385 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-385,-210,-385,-209</points>
<connection>
<GID>856</GID>
<name>IN_0</name></connection>
<intersection>-209 5</intersection></vsegment></shape></wire>
<wire>
<ID>884</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-386,-231,-386,-216</points>
<connection>
<GID>856</GID>
<name>OUT</name></connection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-386,-231,-375.5,-231</points>
<connection>
<GID>817</GID>
<name>K</name></connection>
<intersection>-386 0</intersection></hsegment></shape></wire>
<wire>
<ID>885</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-345,-227.5,-327,-227.5</points>
<connection>
<GID>818</GID>
<name>J</name></connection>
<connection>
<GID>836</GID>
<name>OUT</name></connection>
<intersection>-345 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-345,-227.5,-345,-206.5</points>
<intersection>-227.5 1</intersection>
<intersection>-206.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-345,-206.5,-337.5,-206.5</points>
<intersection>-345 3</intersection>
<intersection>-337.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-337.5,-208,-337.5,-206.5</points>
<connection>
<GID>857</GID>
<name>IN_0</name></connection>
<intersection>-206.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>886</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-338.5,-231.5,-338.5,-214</points>
<connection>
<GID>857</GID>
<name>OUT</name></connection>
<intersection>-231.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-338.5,-231.5,-327,-231.5</points>
<connection>
<GID>818</GID>
<name>K</name></connection>
<intersection>-338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>887</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-592.5,-198,-583.5,-198</points>
<connection>
<GID>867</GID>
<name>IN_1</name></connection>
<connection>
<GID>805</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>888</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-581.5,-198,-581.5,-197</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<intersection>-197 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-575.5,-197,-575.5,-195.5</points>
<connection>
<GID>843</GID>
<name>OUT_0</name></connection>
<intersection>-197 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-581.5,-197,-575.5,-197</points>
<intersection>-581.5 0</intersection>
<intersection>-575.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>889</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-596.5,-247.5,-596.5,-222.5</points>
<intersection>-247.5 1</intersection>
<intersection>-222.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-624,-247.5,-592,-247.5</points>
<connection>
<GID>842</GID>
<name>OUT_0</name></connection>
<connection>
<GID>844</GID>
<name>IN_1</name></connection>
<intersection>-596.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-596.5,-222.5,-591,-222.5</points>
<intersection>-596.5 0</intersection>
<intersection>-591 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-591,-231,-591,-222.5</points>
<connection>
<GID>847</GID>
<name>IN_0</name></connection>
<intersection>-222.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>890</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-610,-245.5,-610,-229.5</points>
<intersection>-245.5 3</intersection>
<intersection>-229.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-624,-229.5,-608.5,-229.5</points>
<connection>
<GID>840</GID>
<name>OUT_0</name></connection>
<intersection>-610 0</intersection>
<intersection>-608.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-610,-245.5,-592,-245.5</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>-610 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-608.5,-230,-608.5,-229.5</points>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<intersection>-229.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-593,-231,-593,-230</points>
<connection>
<GID>847</GID>
<name>IN_1</name></connection>
<intersection>-230 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-604.5,-230,-593,-230</points>
<connection>
<GID>845</GID>
<name>OUT_0</name></connection>
<intersection>-593 0</intersection></hsegment></shape></wire>
<wire>
<ID>892</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-592,-237.5,-586.5,-237.5</points>
<intersection>-592 5</intersection>
<intersection>-586.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-586.5,-237.5,-586.5,-233</points>
<intersection>-237.5 1</intersection>
<intersection>-233 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-592,-237.5,-592,-237</points>
<connection>
<GID>847</GID>
<name>OUT</name></connection>
<intersection>-237.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-586.5,-233,-583,-233</points>
<connection>
<GID>839</GID>
<name>IN_0</name></connection>
<intersection>-586.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>893</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-572.5,-233,-572.5,-216.5</points>
<intersection>-233 1</intersection>
<intersection>-216.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-577,-233,-572.5,-233</points>
<connection>
<GID>839</GID>
<name>OUT_0</name></connection>
<intersection>-572.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-572.5,-216.5,-503,-216.5</points>
<connection>
<GID>820</GID>
<name>IN_0</name></connection>
<intersection>-572.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>894</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-577,-236,-504,-236</points>
<connection>
<GID>821</GID>
<name>IN_1</name></connection>
<connection>
<GID>839</GID>
<name>OUTINV_0</name></connection>
<intersection>-577 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-577,-340.5,-577,-236</points>
<intersection>-340.5 8</intersection>
<intersection>-236 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-577,-340.5,-507,-340.5</points>
<connection>
<GID>858</GID>
<name>IN_3</name></connection>
<intersection>-577 7</intersection></hsegment></shape></wire>
<wire>
<ID>895</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-586,-51,57,-51</points>
<intersection>-586 15</intersection>
<intersection>-578.5 16</intersection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-439.5,57,-51</points>
<intersection>-439.5 3</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-100,-439.5,57,-439.5</points>
<intersection>-100 14</intersection>
<intersection>-84 13</intersection>
<intersection>-70.5 12</intersection>
<intersection>-55.5 11</intersection>
<intersection>-45 10</intersection>
<intersection>-32 9</intersection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-32,-439.5,-32,-428</points>
<connection>
<GID>793</GID>
<name>clock</name></connection>
<intersection>-439.5 3</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-45,-439.5,-45,-428</points>
<connection>
<GID>792</GID>
<name>clock</name></connection>
<intersection>-439.5 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-55.5,-439.5,-55.5,-428</points>
<connection>
<GID>791</GID>
<name>clock</name></connection>
<intersection>-439.5 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-70.5,-439.5,-70.5,-428</points>
<connection>
<GID>790</GID>
<name>clock</name></connection>
<intersection>-439.5 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-84,-439.5,-84,-428</points>
<connection>
<GID>789</GID>
<name>clock</name></connection>
<intersection>-439.5 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-100,-439.5,-100,-427.5</points>
<connection>
<GID>788</GID>
<name>clock</name></connection>
<intersection>-439.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-586,-51,-586,-40.5</points>
<connection>
<GID>910</GID>
<name>CLK</name></connection>
<intersection>-51 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-578.5,-51,-578.5,-40.5</points>
<connection>
<GID>884</GID>
<name>IN_1</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>896</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-330.5,-104,-330.5,-103</points>
<intersection>-104 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-335,-103,-330.5,-103</points>
<connection>
<GID>882</GID>
<name>IN_1</name></connection>
<intersection>-330.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-330.5,-104,-325.5,-104</points>
<connection>
<GID>875</GID>
<name>Q</name></connection>
<intersection>-330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>897</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-561.5,-91.5,-561.5,-87</points>
<intersection>-91.5 1</intersection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-565,-91.5,-561.5,-91.5</points>
<connection>
<GID>889</GID>
<name>IN_1</name></connection>
<intersection>-561.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-561.5,-87,-558,-87</points>
<connection>
<GID>888</GID>
<name>OUT</name></connection>
<intersection>-561.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>898</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-409,-75,-314,-75</points>
<connection>
<GID>871</GID>
<name>OUT_0</name></connection>
<intersection>-314 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-314,-104,-314,-75</points>
<intersection>-104 10</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-319.5,-104,-314,-104</points>
<connection>
<GID>875</GID>
<name>J</name></connection>
<intersection>-314 3</intersection></hsegment></shape></wire>
<wire>
<ID>899</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-571,-104,-341,-104</points>
<connection>
<GID>911</GID>
<name>clear</name></connection>
<connection>
<GID>901</GID>
<name>clear</name></connection>
<connection>
<GID>903</GID>
<name>clear</name></connection>
<connection>
<GID>905</GID>
<name>clear</name></connection>
<connection>
<GID>909</GID>
<name>clear</name></connection>
<connection>
<GID>882</GID>
<name>OUT</name></connection>
<intersection>-571 6</intersection>
<intersection>-434.5 4</intersection>
<intersection>-389 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-389,-104.5,-389,-104</points>
<connection>
<GID>907</GID>
<name>clear</name></connection>
<intersection>-104 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-434.5,-140,-434.5,-104</points>
<intersection>-140 5</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-434.5,-140,-343.5,-140</points>
<intersection>-434.5 4</intersection>
<intersection>-425.5 13</intersection>
<intersection>-409 12</intersection>
<intersection>-394.5 11</intersection>
<intersection>-377.5 10</intersection>
<intersection>-361.5 9</intersection>
<intersection>-343.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-571,-104,-571,-84</points>
<intersection>-104 1</intersection>
<intersection>-84 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-571.5,-84,-571,-84</points>
<connection>
<GID>892</GID>
<name>IN_0</name></connection>
<intersection>-571 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-343.5,-140,-343.5,-139</points>
<connection>
<GID>928</GID>
<name>clear</name></connection>
<intersection>-140 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-361.5,-140,-361.5,-139</points>
<connection>
<GID>927</GID>
<name>clear</name></connection>
<intersection>-140 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-377.5,-140,-377.5,-139</points>
<connection>
<GID>926</GID>
<name>clear</name></connection>
<intersection>-140 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-394.5,-140,-394.5,-139</points>
<connection>
<GID>924</GID>
<name>clear</name></connection>
<intersection>-140 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-409,-140,-409,-139</points>
<connection>
<GID>923</GID>
<name>clear</name></connection>
<intersection>-140 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-425.5,-140,-425.5,-139</points>
<connection>
<GID>921</GID>
<name>clear</name></connection>
<intersection>-140 5</intersection></vsegment></shape></wire>
<wire>
<ID>900</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-565,-93.5,-525,-93.5</points>
<connection>
<GID>889</GID>
<name>IN_0</name></connection>
<intersection>-525 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-525,-95.5,-525,-93.5</points>
<connection>
<GID>886</GID>
<name>OUT</name></connection>
<intersection>-93.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>901</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-583.5,-83,-583.5,-79</points>
<intersection>-83 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-590,-79,-583.5,-79</points>
<connection>
<GID>894</GID>
<name>IN_1</name></connection>
<intersection>-583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-583.5,-83,-577.5,-83</points>
<connection>
<GID>892</GID>
<name>OUT</name></connection>
<intersection>-583.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>902</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-337.5,-100,-337.5,-17</points>
<intersection>-100 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-434,-17,-337.5,-17</points>
<connection>
<GID>879</GID>
<name>IN_0</name></connection>
<intersection>-337.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-337.5,-100,-325.5,-100</points>
<connection>
<GID>875</GID>
<name>nQ</name></connection>
<intersection>-337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>903</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-563,-31,-517.5,-31</points>
<connection>
<GID>893</GID>
<name>clear</name></connection>
<connection>
<GID>891</GID>
<name>clear</name></connection>
<connection>
<GID>890</GID>
<name>clear</name></connection>
<intersection>-563 13</intersection>
<intersection>-517.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-517.5,-32,-517.5,-31</points>
<connection>
<GID>895</GID>
<name>clear</name></connection>
<intersection>-32 5</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-517.5,-32,-436,-32</points>
<connection>
<GID>897</GID>
<name>clear</name></connection>
<connection>
<GID>896</GID>
<name>clear</name></connection>
<intersection>-517.5 4</intersection>
<intersection>-455 12</intersection>
<intersection>-436 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-436,-39,-436,-32</points>
<connection>
<GID>930</GID>
<name>IN_0</name></connection>
<intersection>-32 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-455,-32,-455,-25</points>
<connection>
<GID>898</GID>
<name>OUT</name></connection>
<intersection>-32 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-563,-66,-563,-31</points>
<intersection>-66 14</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-563,-66,-472,-66</points>
<connection>
<GID>936</GID>
<name>clear</name></connection>
<connection>
<GID>935</GID>
<name>clear</name></connection>
<connection>
<GID>934</GID>
<name>clear</name></connection>
<connection>
<GID>933</GID>
<name>clear</name></connection>
<connection>
<GID>932</GID>
<name>clear</name></connection>
<connection>
<GID>931</GID>
<name>clear</name></connection>
<intersection>-563 13</intersection></hsegment></shape></wire>
<wire>
<ID>904</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-467,-12.5,-434,-12.5</points>
<intersection>-467 3</intersection>
<intersection>-434 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-467,-16.5,-467,-12.5</points>
<intersection>-16.5 5</intersection>
<intersection>-12.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-434,-15,-434,-12.5</points>
<connection>
<GID>879</GID>
<name>IN_1</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-468,-16.5,-467,-16.5</points>
<connection>
<GID>925</GID>
<name>OUT</name></connection>
<intersection>-467 3</intersection></hsegment></shape></wire>
<wire>
<ID>905</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-336,-89.5,-336,-87</points>
<intersection>-89.5 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-336,-87,-332,-87</points>
<connection>
<GID>883</GID>
<name>IN_0</name></connection>
<intersection>-336 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-339.5,-89.5,-336,-89.5</points>
<connection>
<GID>920</GID>
<name>OUT</name></connection>
<intersection>-336 0</intersection></hsegment></shape></wire>
<wire>
<ID>906</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-319,-100,-319,-87</points>
<intersection>-100 1</intersection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-319.5,-100,-319,-100</points>
<connection>
<GID>875</GID>
<name>K</name></connection>
<intersection>-319 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-326,-87,-319,-87</points>
<connection>
<GID>883</GID>
<name>OUT_0</name></connection>
<intersection>-319 0</intersection></hsegment></shape></wire>
<wire>
<ID>907</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-582.5,-92.5,-571,-92.5</points>
<connection>
<GID>889</GID>
<name>OUT</name></connection>
<connection>
<GID>902</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-588.5,-91.5,-588.5,-81</points>
<connection>
<GID>902</GID>
<name>OUT</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-590,-81,-588.5,-81</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<intersection>-588.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>909</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-604,-80,-596,-80</points>
<connection>
<GID>894</GID>
<name>OUT</name></connection>
<connection>
<GID>906</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-444.5,-24,-444.5,-16</points>
<intersection>-24 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-449,-24,-444.5,-24</points>
<connection>
<GID>898</GID>
<name>IN_1</name></connection>
<intersection>-444.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-444.5,-16,-440,-16</points>
<connection>
<GID>879</GID>
<name>OUT</name></connection>
<intersection>-444.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-444.5,-108.5,-444.5,-26</points>
<intersection>-108.5 3</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-449,-26,-444.5,-26</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<intersection>-444.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-584,-108.5,-335,-108.5</points>
<connection>
<GID>887</GID>
<name>OUT_0</name></connection>
<intersection>-444.5 0</intersection>
<intersection>-335 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-335,-108.5,-335,-105</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<intersection>-108.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-538,-29,-538,-16.5</points>
<intersection>-29 4</intersection>
<intersection>-25 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-539.5,-16.5,-528.5,-16.5</points>
<connection>
<GID>913</GID>
<name>OUT</name></connection>
<connection>
<GID>916</GID>
<name>IN_0</name></connection>
<intersection>-538 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-538,-25,-536.5,-25</points>
<connection>
<GID>893</GID>
<name>J</name></connection>
<intersection>-538 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-538,-29,-536.5,-29</points>
<connection>
<GID>893</GID>
<name>K</name></connection>
<intersection>-538 0</intersection></hsegment></shape></wire>
<wire>
<ID>913</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-521.5,-29.5,-521.5,-17.5</points>
<intersection>-29.5 4</intersection>
<intersection>-25.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-522.5,-17.5,-513.5,-17.5</points>
<connection>
<GID>916</GID>
<name>OUT</name></connection>
<connection>
<GID>919</GID>
<name>IN_0</name></connection>
<intersection>-521.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-521.5,-25.5,-520.5,-25.5</points>
<connection>
<GID>895</GID>
<name>J</name></connection>
<intersection>-521.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-521.5,-29.5,-520.5,-29.5</points>
<connection>
<GID>895</GID>
<name>K</name></connection>
<intersection>-521.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>914</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-506,-30,-506,-18.5</points>
<intersection>-30 4</intersection>
<intersection>-26 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-507.5,-18.5,-496,-18.5</points>
<connection>
<GID>919</GID>
<name>OUT</name></connection>
<connection>
<GID>922</GID>
<name>IN_0</name></connection>
<intersection>-506 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-506,-26,-504.5,-26</points>
<connection>
<GID>896</GID>
<name>J</name></connection>
<intersection>-506 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-506,-30,-504.5,-30</points>
<connection>
<GID>896</GID>
<name>K</name></connection>
<intersection>-506 0</intersection></hsegment></shape></wire>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-489,-30,-489,-19.5</points>
<intersection>-30 4</intersection>
<intersection>-26 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-490,-19.5,-489,-19.5</points>
<connection>
<GID>922</GID>
<name>OUT</name></connection>
<intersection>-489 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-489,-26,-487.5,-26</points>
<connection>
<GID>897</GID>
<name>J</name></connection>
<intersection>-489 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-489,-30,-487.5,-30</points>
<connection>
<GID>897</GID>
<name>K</name></connection>
<intersection>-489 0</intersection></hsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-560,-25,-552.5,-25</points>
<connection>
<GID>890</GID>
<name>Q</name></connection>
<connection>
<GID>891</GID>
<name>J</name></connection>
<intersection>-559 3</intersection>
<intersection>-556.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-559,-60,-559,-25</points>
<intersection>-60 10</intersection>
<intersection>-44.5 4</intersection>
<intersection>-29 9</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-559,-44.5,-472,-44.5</points>
<connection>
<GID>904</GID>
<name>IN_0</name></connection>
<intersection>-559 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556.5,-25,-556.5,-15.5</points>
<intersection>-25 1</intersection>
<intersection>-15.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-556.5,-15.5,-545.5,-15.5</points>
<connection>
<GID>913</GID>
<name>IN_0</name></connection>
<intersection>-556.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-559,-29,-552.5,-29</points>
<connection>
<GID>891</GID>
<name>K</name></connection>
<intersection>-559 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-559,-60,-557,-60</points>
<connection>
<GID>931</GID>
<name>IN_0</name></connection>
<intersection>-559 3</intersection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-572,-34.5,-317.5,-34.5</points>
<intersection>-572 3</intersection>
<intersection>-556.5 4</intersection>
<intersection>-540.5 32</intersection>
<intersection>-539.5 5</intersection>
<intersection>-526 31</intersection>
<intersection>-523.5 16</intersection>
<intersection>-509 30</intersection>
<intersection>-507 15</intersection>
<intersection>-493 29</intersection>
<intersection>-492 18</intersection>
<intersection>-475 28</intersection>
<intersection>-317.5 35</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-572,-63,-572,-27</points>
<intersection>-63 33</intersection>
<intersection>-39.5 39</intersection>
<intersection>-34.5 1</intersection>
<intersection>-27 13</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-556.5,-34.5,-556.5,-27</points>
<intersection>-34.5 1</intersection>
<intersection>-27 14</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-539.5,-34.5,-539.5,-27</points>
<intersection>-34.5 1</intersection>
<intersection>-27 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-539.5,-27,-536.5,-27</points>
<connection>
<GID>893</GID>
<name>clock</name></connection>
<intersection>-539.5 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-572,-27,-566,-27</points>
<connection>
<GID>890</GID>
<name>clock</name></connection>
<intersection>-572 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-556.5,-27,-552.5,-27</points>
<connection>
<GID>891</GID>
<name>clock</name></connection>
<intersection>-556.5 4</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-507,-34.5,-507,-28</points>
<intersection>-34.5 1</intersection>
<intersection>-28 21</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-523.5,-34.5,-523.5,-27.5</points>
<intersection>-34.5 1</intersection>
<intersection>-27.5 19</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-492,-34.5,-492,-28</points>
<intersection>-34.5 1</intersection>
<intersection>-28 20</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-523.5,-27.5,-520.5,-27.5</points>
<connection>
<GID>895</GID>
<name>clock</name></connection>
<intersection>-523.5 16</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-492,-28,-487.5,-28</points>
<connection>
<GID>897</GID>
<name>clock</name></connection>
<intersection>-492 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-507,-28,-504.5,-28</points>
<connection>
<GID>896</GID>
<name>clock</name></connection>
<intersection>-507 15</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-475,-63,-475,-34.5</points>
<connection>
<GID>936</GID>
<name>clock</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>-493,-63,-493,-34.5</points>
<connection>
<GID>935</GID>
<name>clock</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-509,-63,-509,-34.5</points>
<connection>
<GID>934</GID>
<name>clock</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-526,-63,-526,-34.5</points>
<connection>
<GID>933</GID>
<name>clock</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-540.5,-63,-540.5,-34.5</points>
<connection>
<GID>932</GID>
<name>clock</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-572,-63,-557,-63</points>
<connection>
<GID>931</GID>
<name>clock</name></connection>
<intersection>-572 3</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>-317.5,-102,-317.5,-34.5</points>
<intersection>-102 36</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>-319.5,-102,-317.5,-102</points>
<connection>
<GID>875</GID>
<name>clock</name></connection>
<intersection>-317.5 35</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-572.5,-39.5,-572,-39.5</points>
<connection>
<GID>884</GID>
<name>OUT</name></connection>
<intersection>-572 3</intersection></hsegment></shape></wire>
<wire>
<ID>918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-545.5,-60,-545.5,-17.5</points>
<connection>
<GID>913</GID>
<name>IN_1</name></connection>
<intersection>-60 8</intersection>
<intersection>-43.5 1</intersection>
<intersection>-25 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-545.5,-43.5,-472,-43.5</points>
<connection>
<GID>904</GID>
<name>IN_1</name></connection>
<intersection>-545.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-546.5,-25,-545.5,-25</points>
<connection>
<GID>891</GID>
<name>Q</name></connection>
<intersection>-545.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-545.5,-60,-540.5,-60</points>
<connection>
<GID>932</GID>
<name>IN_0</name></connection>
<intersection>-545.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>919</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-513.5,-41.5,-472,-41.5</points>
<connection>
<GID>904</GID>
<name>IN_3</name></connection>
<intersection>-513.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-513.5,-60,-513.5,-15.5</points>
<connection>
<GID>919</GID>
<name>IN_1</name></connection>
<intersection>-60 9</intersection>
<intersection>-41.5 1</intersection>
<intersection>-25.5 4</intersection>
<intersection>-15.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-514.5,-25.5,-513.5,-25.5</points>
<connection>
<GID>895</GID>
<name>Q</name></connection>
<intersection>-513.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-513.5,-15.5,-474,-15.5</points>
<connection>
<GID>925</GID>
<name>IN_1</name></connection>
<intersection>-513.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-513.5,-60,-509,-60</points>
<connection>
<GID>934</GID>
<name>IN_0</name></connection>
<intersection>-513.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>920</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-529.5,-60,-529.5,-13.5</points>
<intersection>-60 9</intersection>
<intersection>-42.5 4</intersection>
<intersection>-25 3</intersection>
<intersection>-18.5 2</intersection>
<intersection>-13.5 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-529.5,-18.5,-528.5,-18.5</points>
<connection>
<GID>916</GID>
<name>IN_1</name></connection>
<intersection>-529.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-530.5,-25,-529.5,-25</points>
<connection>
<GID>893</GID>
<name>Q</name></connection>
<intersection>-529.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-529.5,-42.5,-472,-42.5</points>
<connection>
<GID>904</GID>
<name>IN_2</name></connection>
<intersection>-529.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-529.5,-13.5,-474,-13.5</points>
<connection>
<GID>925</GID>
<name>IN_0</name></connection>
<intersection>-529.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-529.5,-60,-526,-60</points>
<connection>
<GID>933</GID>
<name>IN_0</name></connection>
<intersection>-529.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-497.5,-60,-497.5,-17.5</points>
<intersection>-60 8</intersection>
<intersection>-40.5 3</intersection>
<intersection>-26 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-498.5,-26,-497.5,-26</points>
<connection>
<GID>896</GID>
<name>Q</name></connection>
<intersection>-497.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-497.5,-17.5,-474,-17.5</points>
<connection>
<GID>925</GID>
<name>IN_2</name></connection>
<intersection>-497.5 0</intersection>
<intersection>-496 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-497.5,-40.5,-472,-40.5</points>
<connection>
<GID>904</GID>
<name>IN_4</name></connection>
<intersection>-497.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-496,-20.5,-496,-17.5</points>
<connection>
<GID>922</GID>
<name>IN_1</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-497.5,-60,-493,-60</points>
<connection>
<GID>935</GID>
<name>IN_0</name></connection>
<intersection>-497.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-479.5,-60,-479.5,-19.5</points>
<intersection>-60 5</intersection>
<intersection>-39.5 2</intersection>
<intersection>-26 1</intersection>
<intersection>-19.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-481.5,-26,-479.5,-26</points>
<connection>
<GID>897</GID>
<name>Q</name></connection>
<intersection>-479.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-479.5,-39.5,-472,-39.5</points>
<connection>
<GID>904</GID>
<name>IN_5</name></connection>
<intersection>-479.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-479.5,-19.5,-474,-19.5</points>
<connection>
<GID>925</GID>
<name>IN_3</name></connection>
<intersection>-479.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-479.5,-60,-475,-60</points>
<connection>
<GID>936</GID>
<name>IN_0</name></connection>
<intersection>-479.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>923</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-549.5,-74.5,-457,-74.5</points>
<connection>
<GID>937</GID>
<name>IN_0</name></connection>
<intersection>-549.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-549.5,-84,-549.5,-60</points>
<intersection>-84 8</intersection>
<intersection>-74.5 1</intersection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-551,-60,-549.5,-60</points>
<connection>
<GID>931</GID>
<name>OUT_0</name></connection>
<intersection>-549.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-551,-84,-549.5,-84</points>
<connection>
<GID>888</GID>
<name>IN_3</name></connection>
<intersection>-549.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>924</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-533,-73.5,-457,-73.5</points>
<connection>
<GID>937</GID>
<name>IN_1</name></connection>
<intersection>-533 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-533,-86,-533,-60</points>
<intersection>-86 8</intersection>
<intersection>-73.5 1</intersection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-534.5,-60,-533,-60</points>
<connection>
<GID>932</GID>
<name>OUT_0</name></connection>
<intersection>-533 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-551,-86,-533,-86</points>
<connection>
<GID>888</GID>
<name>IN_2</name></connection>
<intersection>-533 3</intersection></hsegment></shape></wire>
<wire>
<ID>925</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-519,-72.5,-457,-72.5</points>
<connection>
<GID>937</GID>
<name>IN_2</name></connection>
<intersection>-519 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-519,-88,-519,-60</points>
<intersection>-88 8</intersection>
<intersection>-72.5 1</intersection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-520,-60,-519,-60</points>
<connection>
<GID>933</GID>
<name>OUT_0</name></connection>
<intersection>-519 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-551,-88,-519,-88</points>
<connection>
<GID>888</GID>
<name>IN_1</name></connection>
<intersection>-519 3</intersection></hsegment></shape></wire>
<wire>
<ID>926</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-500.5,-71.5,-457,-71.5</points>
<connection>
<GID>937</GID>
<name>IN_3</name></connection>
<intersection>-500.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-500.5,-90,-500.5,-60</points>
<intersection>-90 8</intersection>
<intersection>-71.5 1</intersection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-503,-60,-500.5,-60</points>
<connection>
<GID>934</GID>
<name>OUT_0</name></connection>
<intersection>-500.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-551,-90,-500.5,-90</points>
<connection>
<GID>888</GID>
<name>IN_0</name></connection>
<intersection>-500.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>927</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-519,-70.5,-457,-70.5</points>
<connection>
<GID>937</GID>
<name>IN_4</name></connection>
<intersection>-519 7</intersection>
<intersection>-486 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-486,-70.5,-486,-60</points>
<intersection>-70.5 1</intersection>
<intersection>-60 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-487,-60,-486,-60</points>
<connection>
<GID>935</GID>
<name>OUT_0</name></connection>
<intersection>-486 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-519,-94.5,-519,-70.5</points>
<connection>
<GID>886</GID>
<name>IN_1</name></connection>
<intersection>-70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-466,-69.5,-457,-69.5</points>
<connection>
<GID>937</GID>
<name>IN_5</name></connection>
<intersection>-466 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-466,-96.5,-466,-60</points>
<intersection>-96.5 8</intersection>
<intersection>-69.5 1</intersection>
<intersection>-60 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-469,-60,-466,-60</points>
<connection>
<GID>936</GID>
<name>OUT_0</name></connection>
<intersection>-466 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-519,-96.5,-466,-96.5</points>
<connection>
<GID>886</GID>
<name>IN_0</name></connection>
<intersection>-466 5</intersection></hsegment></shape></wire>
<wire>
<ID>929</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-409.5,-102,-409.5,-89.5</points>
<intersection>-102 4</intersection>
<intersection>-98 2</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-411,-89.5,-400,-89.5</points>
<connection>
<GID>914</GID>
<name>OUT</name></connection>
<connection>
<GID>915</GID>
<name>IN_0</name></connection>
<intersection>-409.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-409.5,-98,-408,-98</points>
<connection>
<GID>905</GID>
<name>J</name></connection>
<intersection>-409.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-409.5,-102,-408,-102</points>
<connection>
<GID>905</GID>
<name>K</name></connection>
<intersection>-409.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-393,-102.5,-393,-90.5</points>
<intersection>-102.5 4</intersection>
<intersection>-98.5 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-394,-90.5,-385,-90.5</points>
<connection>
<GID>915</GID>
<name>OUT</name></connection>
<connection>
<GID>917</GID>
<name>IN_0</name></connection>
<intersection>-393 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-393,-98.5,-392,-98.5</points>
<connection>
<GID>907</GID>
<name>J</name></connection>
<intersection>-393 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-393,-102.5,-392,-102.5</points>
<connection>
<GID>907</GID>
<name>K</name></connection>
<intersection>-393 0</intersection></hsegment></shape></wire>
<wire>
<ID>931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-377.5,-102,-377.5,-91.5</points>
<intersection>-102 4</intersection>
<intersection>-98 2</intersection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-379,-91.5,-367.5,-91.5</points>
<connection>
<GID>917</GID>
<name>OUT</name></connection>
<connection>
<GID>918</GID>
<name>IN_0</name></connection>
<intersection>-377.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-377.5,-98,-376,-98</points>
<connection>
<GID>909</GID>
<name>J</name></connection>
<intersection>-377.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-377.5,-102,-376,-102</points>
<connection>
<GID>909</GID>
<name>K</name></connection>
<intersection>-377.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-360.5,-102,-360.5,-92.5</points>
<intersection>-102 4</intersection>
<intersection>-98 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-361.5,-92.5,-360.5,-92.5</points>
<connection>
<GID>918</GID>
<name>OUT</name></connection>
<intersection>-360.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-360.5,-98,-359,-98</points>
<connection>
<GID>911</GID>
<name>J</name></connection>
<intersection>-360.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-360.5,-102,-359,-102</points>
<connection>
<GID>911</GID>
<name>K</name></connection>
<intersection>-360.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-431.5,-98,-424,-98</points>
<connection>
<GID>901</GID>
<name>Q</name></connection>
<connection>
<GID>903</GID>
<name>J</name></connection>
<intersection>-430.5 3</intersection>
<intersection>-428 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-430.5,-133,-430.5,-98</points>
<intersection>-133 10</intersection>
<intersection>-117.5 4</intersection>
<intersection>-102 9</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-430.5,-117.5,-349,-117.5</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<intersection>-430.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-428,-98,-428,-88.5</points>
<intersection>-98 1</intersection>
<intersection>-88.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-428,-88.5,-417,-88.5</points>
<connection>
<GID>914</GID>
<name>IN_0</name></connection>
<intersection>-428 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-430.5,-102,-424,-102</points>
<connection>
<GID>903</GID>
<name>K</name></connection>
<intersection>-430.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-430.5,-133,-428.5,-133</points>
<connection>
<GID>921</GID>
<name>IN_0</name></connection>
<intersection>-430.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-417,-133,-417,-90.5</points>
<connection>
<GID>914</GID>
<name>IN_1</name></connection>
<intersection>-133 8</intersection>
<intersection>-116.5 1</intersection>
<intersection>-98 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-417,-116.5,-349,-116.5</points>
<connection>
<GID>912</GID>
<name>IN_1</name></connection>
<intersection>-417 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-418,-98,-417,-98</points>
<connection>
<GID>903</GID>
<name>Q</name></connection>
<intersection>-417 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-417,-133,-412,-133</points>
<connection>
<GID>923</GID>
<name>IN_0</name></connection>
<intersection>-417 0</intersection></hsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-385,-114.5,-349,-114.5</points>
<connection>
<GID>912</GID>
<name>IN_3</name></connection>
<intersection>-385 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-385,-133,-385,-88.5</points>
<connection>
<GID>917</GID>
<name>IN_1</name></connection>
<intersection>-133 9</intersection>
<intersection>-114.5 1</intersection>
<intersection>-98.5 4</intersection>
<intersection>-88.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-386,-98.5,-385,-98.5</points>
<connection>
<GID>907</GID>
<name>Q</name></connection>
<intersection>-385 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-385,-88.5,-345.5,-88.5</points>
<connection>
<GID>920</GID>
<name>IN_1</name></connection>
<intersection>-385 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-385,-133,-380.5,-133</points>
<connection>
<GID>926</GID>
<name>IN_0</name></connection>
<intersection>-385 3</intersection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-401,-133,-401,-86.5</points>
<intersection>-133 9</intersection>
<intersection>-115.5 4</intersection>
<intersection>-98 3</intersection>
<intersection>-91.5 2</intersection>
<intersection>-86.5 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-401,-91.5,-400,-91.5</points>
<connection>
<GID>915</GID>
<name>IN_1</name></connection>
<intersection>-401 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-402,-98,-401,-98</points>
<connection>
<GID>905</GID>
<name>Q</name></connection>
<intersection>-401 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-401,-115.5,-349,-115.5</points>
<connection>
<GID>912</GID>
<name>IN_2</name></connection>
<intersection>-401 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-401,-86.5,-345.5,-86.5</points>
<connection>
<GID>920</GID>
<name>IN_0</name></connection>
<intersection>-401 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-401,-133,-397.5,-133</points>
<connection>
<GID>924</GID>
<name>IN_0</name></connection>
<intersection>-401 0</intersection></hsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-369,-133,-369,-90.5</points>
<intersection>-133 8</intersection>
<intersection>-113.5 3</intersection>
<intersection>-98 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-370,-98,-369,-98</points>
<connection>
<GID>909</GID>
<name>Q</name></connection>
<intersection>-369 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-369,-90.5,-345.5,-90.5</points>
<connection>
<GID>920</GID>
<name>IN_2</name></connection>
<intersection>-369 0</intersection>
<intersection>-367.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-369,-113.5,-349,-113.5</points>
<connection>
<GID>912</GID>
<name>IN_4</name></connection>
<intersection>-369 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-367.5,-93.5,-367.5,-90.5</points>
<connection>
<GID>918</GID>
<name>IN_1</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-369,-133,-364.5,-133</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<intersection>-369 0</intersection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-351,-133,-351,-92.5</points>
<intersection>-133 5</intersection>
<intersection>-112.5 2</intersection>
<intersection>-98 1</intersection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-353,-98,-351,-98</points>
<connection>
<GID>911</GID>
<name>Q</name></connection>
<intersection>-351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-351,-112.5,-349,-112.5</points>
<connection>
<GID>912</GID>
<name>IN_5</name></connection>
<intersection>-351 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-351,-92.5,-345.5,-92.5</points>
<connection>
<GID>920</GID>
<name>IN_3</name></connection>
<intersection>-351 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-351,-133,-346.5,-133</points>
<connection>
<GID>928</GID>
<name>IN_0</name></connection>
<intersection>-351 0</intersection></hsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-421,-185,-100,-185</points>
<intersection>-421 3</intersection>
<intersection>-100 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-421,-185,-421,-133</points>
<intersection>-185 1</intersection>
<intersection>-147.5 7</intersection>
<intersection>-133 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-422.5,-133,-421,-133</points>
<connection>
<GID>921</GID>
<name>OUT_0</name></connection>
<intersection>-421 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-100,-415,-100,-185</points>
<connection>
<GID>940</GID>
<name>IN_0</name></connection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-421,-147.5,-328.5,-147.5</points>
<connection>
<GID>929</GID>
<name>IN_0</name></connection>
<intersection>-421 3</intersection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-404.5,-180.5,-86.5,-180.5</points>
<intersection>-404.5 3</intersection>
<intersection>-86.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-404.5,-180.5,-404.5,-133</points>
<intersection>-180.5 1</intersection>
<intersection>-146.5 7</intersection>
<intersection>-133 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-406,-133,-404.5,-133</points>
<connection>
<GID>923</GID>
<name>OUT_0</name></connection>
<intersection>-404.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-86.5,-415,-86.5,-180.5</points>
<connection>
<GID>942</GID>
<name>IN_0</name></connection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-404.5,-146.5,-328.5,-146.5</points>
<connection>
<GID>929</GID>
<name>IN_1</name></connection>
<intersection>-404.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-390.5,-176,-73.5,-176</points>
<intersection>-390.5 3</intersection>
<intersection>-73.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-390.5,-176,-390.5,-133</points>
<intersection>-176 1</intersection>
<intersection>-145.5 7</intersection>
<intersection>-133 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-391.5,-133,-390.5,-133</points>
<connection>
<GID>924</GID>
<name>OUT_0</name></connection>
<intersection>-390.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-73.5,-415,-73.5,-176</points>
<connection>
<GID>943</GID>
<name>IN_0</name></connection>
<intersection>-176 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-390.5,-145.5,-328.5,-145.5</points>
<connection>
<GID>929</GID>
<name>IN_2</name></connection>
<intersection>-390.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-372,-171.5,-60.5,-171.5</points>
<intersection>-372 3</intersection>
<intersection>-60.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-372,-171.5,-372,-133</points>
<intersection>-171.5 1</intersection>
<intersection>-144.5 7</intersection>
<intersection>-133 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-374.5,-133,-372,-133</points>
<connection>
<GID>926</GID>
<name>OUT_0</name></connection>
<intersection>-372 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-60.5,-415,-60.5,-171.5</points>
<connection>
<GID>945</GID>
<name>IN_0</name></connection>
<intersection>-171.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-372,-144.5,-328.5,-144.5</points>
<connection>
<GID>929</GID>
<name>IN_3</name></connection>
<intersection>-372 3</intersection></hsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-357,-168.5,-48,-168.5</points>
<intersection>-357 3</intersection>
<intersection>-48 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-357,-168.5,-357,-133</points>
<intersection>-168.5 1</intersection>
<intersection>-143.5 7</intersection>
<intersection>-133 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-358.5,-133,-357,-133</points>
<connection>
<GID>927</GID>
<name>OUT_0</name></connection>
<intersection>-357 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-48,-415.5,-48,-168.5</points>
<connection>
<GID>947</GID>
<name>IN_0</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-357,-143.5,-328.5,-143.5</points>
<connection>
<GID>929</GID>
<name>IN_4</name></connection>
<intersection>-357 3</intersection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-334.5,-163.5,-334.5,-133</points>
<intersection>-163.5 5</intersection>
<intersection>-142.5 8</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-340.5,-133,-334.5,-133</points>
<connection>
<GID>928</GID>
<name>OUT_0</name></connection>
<intersection>-334.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-334.5,-163.5,-35.5,-163.5</points>
<intersection>-334.5 0</intersection>
<intersection>-35.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-35.5,-415.5,-35.5,-163.5</points>
<connection>
<GID>948</GID>
<name>IN_0</name></connection>
<intersection>-163.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-334.5,-142.5,-328.5,-142.5</points>
<connection>
<GID>929</GID>
<name>IN_5</name></connection>
<intersection>-334.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-441,-102,-441,-75</points>
<intersection>-102 4</intersection>
<intersection>-98 17</intersection>
<intersection>-75 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-580,-102,-437.5,-102</points>
<connection>
<GID>901</GID>
<name>K</name></connection>
<intersection>-580 11</intersection>
<intersection>-441 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-441,-75,-415,-75</points>
<connection>
<GID>871</GID>
<name>IN_0</name></connection>
<intersection>-441 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-580,-25,-566,-25</points>
<connection>
<GID>890</GID>
<name>J</name></connection>
<intersection>-580 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-580,-102,-580,-25</points>
<intersection>-102 4</intersection>
<intersection>-90.5 22</intersection>
<intersection>-77.5 23</intersection>
<intersection>-38.5 21</intersection>
<intersection>-31 28</intersection>
<intersection>-29 14</intersection>
<intersection>-25 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-580,-29,-566,-29</points>
<connection>
<GID>890</GID>
<name>K</name></connection>
<intersection>-580 11</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-441,-98,-437.5,-98</points>
<connection>
<GID>901</GID>
<name>J</name></connection>
<intersection>-441 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-580,-38.5,-578.5,-38.5</points>
<connection>
<GID>884</GID>
<name>IN_0</name></connection>
<intersection>-580 11</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-582.5,-90.5,-580,-90.5</points>
<connection>
<GID>902</GID>
<name>IN_1</name></connection>
<intersection>-580 11</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-580,-77.5,-571.5,-77.5</points>
<intersection>-580 11</intersection>
<intersection>-571.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-571.5,-82,-571.5,-77.5</points>
<connection>
<GID>892</GID>
<name>IN_1</name></connection>
<intersection>-77.5 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-586.5,-31,-580,-31</points>
<connection>
<GID>938</GID>
<name>OUT</name></connection>
<intersection>-580 11</intersection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-438.5,-136,-438.5,-45</points>
<intersection>-136 8</intersection>
<intersection>-100 1</intersection>
<intersection>-45 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-438.5,-100,-359,-100</points>
<connection>
<GID>901</GID>
<name>clock</name></connection>
<connection>
<GID>903</GID>
<name>clock</name></connection>
<connection>
<GID>905</GID>
<name>clock</name></connection>
<connection>
<GID>909</GID>
<name>clock</name></connection>
<connection>
<GID>911</GID>
<name>clock</name></connection>
<intersection>-438.5 0</intersection>
<intersection>-392 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-392,-100.5,-392,-100</points>
<connection>
<GID>907</GID>
<name>clock</name></connection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-438.5,-136,-346.5,-136</points>
<connection>
<GID>921</GID>
<name>clock</name></connection>
<connection>
<GID>923</GID>
<name>clock</name></connection>
<connection>
<GID>924</GID>
<name>clock</name></connection>
<connection>
<GID>926</GID>
<name>clock</name></connection>
<connection>
<GID>927</GID>
<name>clock</name></connection>
<connection>
<GID>928</GID>
<name>clock</name></connection>
<intersection>-438.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-438.5,-45,-436,-45</points>
<connection>
<GID>930</GID>
<name>OUT_0</name></connection>
<intersection>-438.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>181.017,265.324,1405.02,-339.676</PageViewport>
<gate>
<ID>950</ID>
<type>CC_PULSE</type>
<position>323,-96</position>
<output>
<ID>OUT_0</ID>1053 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>951</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>670,-147.5</position>
<input>
<ID>IN_0</ID>1005 </input>
<input>
<ID>IN_1</ID>1023 </input>
<input>
<ID>IN_2</ID>1024 </input>
<input>
<ID>IN_3</ID>1025 </input>
<input>
<ID>IN_4</ID>1026 </input>
<input>
<ID>IN_5</ID>1027 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>952</ID>
<type>CC_PULSE</type>
<position>324,-114</position>
<output>
<ID>OUT_0</ID>1052 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>953</ID>
<type>EE_VDD</type>
<position>374.5,-61</position>
<output>
<ID>OUT_0</ID>1051 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>954</ID>
<type>AE_OR2</type>
<position>361,-113</position>
<input>
<ID>IN_0</ID>1053 </input>
<input>
<ID>IN_1</ID>1052 </input>
<output>
<ID>OUT</ID>1021 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>955</ID>
<type>AE_DFF_LOW</type>
<position>869,-293.5</position>
<input>
<ID>IN_0</ID>969 </input>
<output>
<ID>OUT_0</ID>975 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>956</ID>
<type>AE_SMALL_INVERTER</type>
<position>343.5,-96.5</position>
<input>
<ID>IN_0</ID>1053 </input>
<output>
<ID>OUT_0</ID>1054 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>957</ID>
<type>AA_AND2</type>
<position>467.5,-188</position>
<input>
<ID>IN_0</ID>1032 </input>
<input>
<ID>IN_1</ID>1031 </input>
<output>
<ID>OUT</ID>1033 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>958</ID>
<type>AI_XOR2</type>
<position>358,-100.5</position>
<input>
<ID>IN_0</ID>1052 </input>
<input>
<ID>IN_1</ID>1054 </input>
<output>
<ID>OUT</ID>1055 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>959</ID>
<type>AA_LABEL</type>
<position>328,-90</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>960</ID>
<type>AA_AND2</type>
<position>541.5,-174.5</position>
<input>
<ID>IN_0</ID>1034 </input>
<input>
<ID>IN_1</ID>1035 </input>
<output>
<ID>OUT</ID>1036 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>961</ID>
<type>AA_LABEL</type>
<position>327,-119</position>
<gparam>LABEL_TEXT Decrement</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>962</ID>
<type>AA_AND2</type>
<position>604.5,-173</position>
<input>
<ID>IN_0</ID>1037 </input>
<input>
<ID>IN_1</ID>1038 </input>
<output>
<ID>OUT</ID>1039 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>963</ID>
<type>AI_XOR2</type>
<position>418,-82</position>
<input>
<ID>IN_0</ID>1028 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1030 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>964</ID>
<type>AE_DFF_LOW</type>
<position>882.5,-293.5</position>
<input>
<ID>IN_0</ID>970 </input>
<output>
<ID>OUT_0</ID>976 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>965</ID>
<type>AI_XOR2</type>
<position>469,-79.5</position>
<input>
<ID>IN_0</ID>1040 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1041 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>966</ID>
<type>AI_XOR2</type>
<position>505.5,-79</position>
<input>
<ID>IN_0</ID>1043 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1042 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>967</ID>
<type>AI_XOR2</type>
<position>534,-79.5</position>
<input>
<ID>IN_0</ID>1044 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1045 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>968</ID>
<type>AI_XOR2</type>
<position>564,-79.5</position>
<input>
<ID>IN_0</ID>1046 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1047 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>969</ID>
<type>AI_XOR2</type>
<position>611.5,-77.5</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1049 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>970</ID>
<type>AA_AND4</type>
<position>446,-210</position>
<input>
<ID>IN_0</ID>1039 </input>
<input>
<ID>IN_1</ID>1036 </input>
<input>
<ID>IN_2</ID>1033 </input>
<input>
<ID>IN_3</ID>1057 </input>
<output>
<ID>OUT</ID>1029 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>971</ID>
<type>AE_DFF_LOW</type>
<position>897.5,-293.5</position>
<input>
<ID>IN_0</ID>971 </input>
<output>
<ID>OUT_0</ID>977 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>972</ID>
<type>AA_INVERTER</type>
<position>461.5,-165</position>
<input>
<ID>IN_0</ID>1000 </input>
<output>
<ID>OUT_0</ID>1031 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>973</ID>
<type>AA_INVERTER</type>
<position>474,-166</position>
<input>
<ID>IN_0</ID>1004 </input>
<output>
<ID>OUT_0</ID>1032 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>974</ID>
<type>AA_INVERTER</type>
<position>538,-165</position>
<input>
<ID>IN_0</ID>1009 </input>
<output>
<ID>OUT_0</ID>1035 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>975</ID>
<type>AA_INVERTER</type>
<position>545,-165</position>
<input>
<ID>IN_0</ID>1013 </input>
<output>
<ID>OUT_0</ID>1034 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>976</ID>
<type>AE_DFF_LOW</type>
<position>908,-293.5</position>
<input>
<ID>IN_0</ID>972 </input>
<output>
<ID>OUT_0</ID>978 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>977</ID>
<type>AA_INVERTER</type>
<position>602.5,-164.5</position>
<input>
<ID>IN_0</ID>1017 </input>
<output>
<ID>OUT_0</ID>1038 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>978</ID>
<type>AA_INVERTER</type>
<position>608,-164</position>
<input>
<ID>IN_0</ID>1022 </input>
<output>
<ID>OUT_0</ID>1037 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>979</ID>
<type>AA_LABEL</type>
<position>670,-157.5</position>
<gparam>LABEL_TEXT Actual Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>980</ID>
<type>AA_AND2</type>
<position>367.5,-67.5</position>
<input>
<ID>IN_0</ID>1051 </input>
<input>
<ID>IN_1</ID>1050 </input>
<output>
<ID>OUT</ID>1028 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>981</ID>
<type>AA_LABEL</type>
<position>496.5,-58</position>
<gparam>LABEL_TEXT Setting Mode</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>982</ID>
<type>AE_DFF_LOW</type>
<position>921,-293.5</position>
<input>
<ID>IN_0</ID>973 </input>
<output>
<ID>OUT_0</ID>979 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>983</ID>
<type>AA_LABEL</type>
<position>361.5,-54.5</position>
<gparam>LABEL_TEXT On/Off- Settings/Cycle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>984</ID>
<type>AA_INVERTER</type>
<position>538,58.5</position>
<input>
<ID>IN_0</ID>1108 </input>
<output>
<ID>OUT_0</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>985</ID>
<type>AA_LABEL</type>
<position>348,134</position>
<gparam>LABEL_TEXT Water Button</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>986</ID>
<type>AE_SMALL_INVERTER</type>
<position>860,-301</position>
<input>
<ID>IN_0</ID>974 </input>
<output>
<ID>OUT_0</ID>980 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>987</ID>
<type>AA_LABEL</type>
<position>498.5,93</position>
<gparam>LABEL_TEXT Buffer Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>988</ID>
<type>AA_LABEL</type>
<position>440.5,144.5</position>
<gparam>LABEL_TEXT Seconds Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>989</ID>
<type>AE_SMALL_INVERTER</type>
<position>875,-301</position>
<input>
<ID>IN_0</ID>975 </input>
<output>
<ID>OUT_0</ID>981 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>990</ID>
<type>BE_JKFF_LOW_NT</type>
<position>627.5,31.5</position>
<input>
<ID>J</ID>1061 </input>
<input>
<ID>K</ID>1069 </input>
<output>
<ID>Q</ID>1059 </output>
<input>
<ID>clock</ID>1080 </input>
<output>
<ID>nQ</ID>1065 </output>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>991</ID>
<type>AA_LABEL</type>
<position>497,71.5</position>
<gparam>LABEL_TEXT Actual Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>992</ID>
<type>AE_SMALL_INVERTER</type>
<position>890,-301</position>
<input>
<ID>IN_0</ID>976 </input>
<output>
<ID>OUT_0</ID>982 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>993</ID>
<type>AA_LABEL</type>
<position>571,53</position>
<gparam>LABEL_TEXT Minutes Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>994</ID>
<type>AE_SMALL_INVERTER</type>
<position>901.5,-300.5</position>
<input>
<ID>IN_0</ID>977 </input>
<output>
<ID>OUT_0</ID>983 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>995</ID>
<type>AA_LABEL</type>
<position>634,17.5</position>
<gparam>LABEL_TEXT Buffer Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>996</ID>
<type>AE_SMALL_INVERTER</type>
<position>914.5,-301</position>
<input>
<ID>IN_0</ID>978 </input>
<output>
<ID>OUT_0</ID>984 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>997</ID>
<type>AI_XOR2</type>
<position>513,117.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<input>
<ID>IN_1</ID>1067 </input>
<output>
<ID>OUT</ID>1073 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>998</ID>
<type>AA_LABEL</type>
<position>517.5,127.5</position>
<gparam>LABEL_TEXT Both on seconds counter stop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>999</ID>
<type>AE_SMALL_INVERTER</type>
<position>927.5,-300.5</position>
<input>
<ID>IN_0</ID>979 </input>
<output>
<ID>OUT_0</ID>985 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1000</ID>
<type>AA_LABEL</type>
<position>643.5,-11.5</position>
<gparam>LABEL_TEXT Actual Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1001</ID>
<type>AI_XOR2</type>
<position>612,29.5</position>
<input>
<ID>IN_0</ID>1074 </input>
<input>
<ID>IN_1</ID>1059 </input>
<output>
<ID>OUT</ID>1062 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1002</ID>
<type>AA_INVERTER</type>
<position>621,46.5</position>
<input>
<ID>IN_0</ID>1068 </input>
<output>
<ID>OUT_0</ID>1069 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1003</ID>
<type>AA_AND2</type>
<position>374.5,94</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1058 </input>
<output>
<ID>OUT</ID>1080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1004</ID>
<type>AA_LABEL</type>
<position>363.5,20</position>
<gparam>LABEL_TEXT Abort</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1005</ID>
<type>AE_OR2</type>
<position>428,38</position>
<input>
<ID>IN_0</ID>1091 </input>
<input>
<ID>IN_1</ID>1090 </input>
<output>
<ID>OUT</ID>1063 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1006</ID>
<type>AA_TOGGLE</type>
<position>364,25</position>
<output>
<ID>OUT_0</ID>1074 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1007</ID>
<type>AE_OR4</type>
<position>396,46.5</position>
<input>
<ID>IN_0</ID>1089 </input>
<input>
<ID>IN_1</ID>1088 </input>
<input>
<ID>IN_2</ID>1087 </input>
<input>
<ID>IN_3</ID>1086 </input>
<output>
<ID>OUT</ID>1060 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1008</ID>
<type>AE_OR2</type>
<position>382,41</position>
<input>
<ID>IN_0</ID>1063 </input>
<input>
<ID>IN_1</ID>1060 </input>
<output>
<ID>OUT</ID>1070 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1009</ID>
<type>BE_JKFF_LOW_NT</type>
<position>387,106.5</position>
<input>
<ID>J</ID>1108 </input>
<input>
<ID>K</ID>1108 </input>
<output>
<ID>Q</ID>1079 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1010</ID>
<type>BE_JKFF_LOW_NT</type>
<position>400.5,106.5</position>
<input>
<ID>J</ID>1079 </input>
<input>
<ID>K</ID>1079 </input>
<output>
<ID>Q</ID>1081 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1011</ID>
<type>AA_AND2</type>
<position>375.5,50.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<input>
<ID>IN_1</ID>1108 </input>
<output>
<ID>OUT</ID>1064 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1012</ID>
<type>BE_JKFF_LOW_NT</type>
<position>416.5,106.5</position>
<input>
<ID>J</ID>1075 </input>
<input>
<ID>K</ID>1075 </input>
<output>
<ID>Q</ID>1083 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1013</ID>
<type>AA_TOGGLE</type>
<position>729,-185</position>
<output>
<ID>OUT_0</ID>967 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1014</ID>
<type>AE_OR2</type>
<position>357,53.5</position>
<input>
<ID>IN_0</ID>1071 </input>
<input>
<ID>IN_1</ID>1064 </input>
<output>
<ID>OUT</ID>1072 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1015</ID>
<type>BE_JKFF_LOW_NT</type>
<position>432.5,106</position>
<input>
<ID>J</ID>1076 </input>
<input>
<ID>K</ID>1076 </input>
<output>
<ID>Q</ID>1082 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1016</ID>
<type>AA_AND4</type>
<position>878,-317.5</position>
<input>
<ID>IN_0</ID>983 </input>
<input>
<ID>IN_1</ID>982 </input>
<input>
<ID>IN_2</ID>981 </input>
<input>
<ID>IN_3</ID>980 </input>
<output>
<ID>OUT</ID>986 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1017</ID>
<type>BE_JKFF_LOW_NT</type>
<position>448.5,105.5</position>
<input>
<ID>J</ID>1077 </input>
<input>
<ID>K</ID>1077 </input>
<output>
<ID>Q</ID>1084 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1018</ID>
<type>BE_JKFF_LOW_NT</type>
<position>465.5,105.5</position>
<input>
<ID>J</ID>1078 </input>
<input>
<ID>K</ID>1078 </input>
<output>
<ID>Q</ID>1085 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1019</ID>
<type>AI_XOR2</type>
<position>498,108.5</position>
<input>
<ID>IN_0</ID>1074 </input>
<input>
<ID>IN_1</ID>1073 </input>
<output>
<ID>OUT</ID>1066 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1020</ID>
<type>AA_TOGGLE</type>
<position>356.5,126.5</position>
<output>
<ID>OUT_0</ID>988 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1021</ID>
<type>AA_LABEL</type>
<position>343.5,60.5</position>
<gparam>LABEL_TEXT Water On/Off</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1022</ID>
<type>BE_JKFF_LOW_NT</type>
<position>515.5,33.5</position>
<input>
<ID>J</ID>1108 </input>
<input>
<ID>K</ID>1108 </input>
<output>
<ID>Q</ID>1096 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1023</ID>
<type>AA_AND2</type>
<position>364.5,42</position>
<input>
<ID>IN_0</ID>1070 </input>
<input>
<ID>IN_1</ID>1108 </input>
<output>
<ID>OUT</ID>1071 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1024</ID>
<type>BE_JKFF_LOW_NT</type>
<position>529,33.5</position>
<input>
<ID>J</ID>1096 </input>
<input>
<ID>K</ID>1096 </input>
<output>
<ID>Q</ID>1097 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1025</ID>
<type>AE_DFF_LOW</type>
<position>870,-408.5</position>
<input>
<ID>IN_0</ID>948 </input>
<output>
<ID>OUT_0</ID>954 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1026</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>483,92</position>
<input>
<ID>IN_0</ID>1079 </input>
<input>
<ID>IN_1</ID>1081 </input>
<input>
<ID>IN_2</ID>1083 </input>
<input>
<ID>IN_3</ID>1082 </input>
<input>
<ID>IN_4</ID>1084 </input>
<input>
<ID>IN_5</ID>1085 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1027</ID>
<type>BE_JKFF_LOW_NT</type>
<position>545,33.5</position>
<input>
<ID>J</ID>1092 </input>
<input>
<ID>K</ID>1092 </input>
<output>
<ID>Q</ID>1099 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1028</ID>
<type>AA_AND2</type>
<position>914.5,-316.5</position>
<input>
<ID>IN_0</ID>985 </input>
<input>
<ID>IN_1</ID>984 </input>
<output>
<ID>OUT</ID>987 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1029</ID>
<type>GA_LED</type>
<position>345,53.5</position>
<input>
<ID>N_in1</ID>1072 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1030</ID>
<type>BE_JKFF_LOW_NT</type>
<position>561,33</position>
<input>
<ID>J</ID>1093 </input>
<input>
<ID>K</ID>1093 </input>
<output>
<ID>Q</ID>1098 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1031</ID>
<type>AA_AND2</type>
<position>893.5,-329.5</position>
<input>
<ID>IN_0</ID>987 </input>
<input>
<ID>IN_1</ID>986 </input>
<output>
<ID>OUT</ID>990 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1032</ID>
<type>AA_LABEL</type>
<position>395.5,35.5</position>
<gparam>LABEL_TEXT Output of Flip-flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1033</ID>
<type>BE_JKFF_LOW_NT</type>
<position>577,33.5</position>
<input>
<ID>J</ID>1094 </input>
<input>
<ID>K</ID>1094 </input>
<output>
<ID>Q</ID>1100 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1034</ID>
<type>BB_CLOCK</type>
<position>360,93</position>
<output>
<ID>CLK</ID>1058 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 3</lparam></gate>
<gate>
<ID>1035</ID>
<type>BE_JKFF_LOW_NT</type>
<position>594,33.5</position>
<input>
<ID>J</ID>1095 </input>
<input>
<ID>K</ID>1095 </input>
<output>
<ID>Q</ID>1101 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1036</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>606,19</position>
<input>
<ID>IN_0</ID>1096 </input>
<input>
<ID>IN_1</ID>1097 </input>
<input>
<ID>IN_2</ID>1099 </input>
<input>
<ID>IN_3</ID>1098 </input>
<input>
<ID>IN_4</ID>1100 </input>
<input>
<ID>IN_5</ID>1101 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1037</ID>
<type>AA_AND2</type>
<position>407.5,117</position>
<input>
<ID>IN_0</ID>1079 </input>
<input>
<ID>IN_1</ID>1081 </input>
<output>
<ID>OUT</ID>1075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1038</ID>
<type>AI_XOR2</type>
<position>369,119</position>
<input>
<ID>IN_0</ID>990 </input>
<input>
<ID>IN_1</ID>988 </input>
<output>
<ID>OUT</ID>989 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1039</ID>
<type>AE_DFF_LOW</type>
<position>883.5,-408.5</position>
<input>
<ID>IN_0</ID>949 </input>
<output>
<ID>OUT_0</ID>955 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1040</ID>
<type>AA_AND2</type>
<position>536,44</position>
<input>
<ID>IN_0</ID>1096 </input>
<input>
<ID>IN_1</ID>1097 </input>
<output>
<ID>OUT</ID>1092 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1041</ID>
<type>AA_AND2</type>
<position>553,43</position>
<input>
<ID>IN_0</ID>1092 </input>
<input>
<ID>IN_1</ID>1099 </input>
<output>
<ID>OUT</ID>1093 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1042</ID>
<type>AA_AND2</type>
<position>424.5,116</position>
<input>
<ID>IN_0</ID>1075 </input>
<input>
<ID>IN_1</ID>1083 </input>
<output>
<ID>OUT</ID>1076 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1043</ID>
<type>AA_AND2</type>
<position>568,42</position>
<input>
<ID>IN_0</ID>1093 </input>
<input>
<ID>IN_1</ID>1098 </input>
<output>
<ID>OUT</ID>1094 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1044</ID>
<type>AE_DFF_LOW</type>
<position>898.5,-408.5</position>
<input>
<ID>IN_0</ID>950 </input>
<output>
<ID>OUT_0</ID>956 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1045</ID>
<type>AA_AND2</type>
<position>585.5,41</position>
<input>
<ID>IN_0</ID>1094 </input>
<input>
<ID>IN_1</ID>1100 </input>
<output>
<ID>OUT</ID>1095 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1046</ID>
<type>AA_AND2</type>
<position>439.5,115</position>
<input>
<ID>IN_0</ID>1076 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1077 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1047</ID>
<type>BA_NAND4</type>
<position>607.5,44</position>
<input>
<ID>IN_0</ID>1099 </input>
<input>
<ID>IN_1</ID>1098 </input>
<input>
<ID>IN_2</ID>1100 </input>
<input>
<ID>IN_3</ID>1101 </input>
<output>
<ID>OUT</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1048</ID>
<type>AE_DFF_LOW</type>
<position>524.5,-1.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<output>
<ID>OUT_0</ID>1102 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1049</ID>
<type>AA_AND2</type>
<position>457,114</position>
<input>
<ID>IN_0</ID>1077 </input>
<input>
<ID>IN_1</ID>1084 </input>
<output>
<ID>OUT</ID>1078 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1050</ID>
<type>AE_DFF_LOW</type>
<position>909,-408.5</position>
<input>
<ID>IN_0</ID>951 </input>
<output>
<ID>OUT_0</ID>957 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1051</ID>
<type>AE_DFF_LOW</type>
<position>541,-1.5</position>
<input>
<ID>IN_0</ID>1097 </input>
<output>
<ID>OUT_0</ID>1103 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1052</ID>
<type>AE_DFF_LOW</type>
<position>922,-408.5</position>
<input>
<ID>IN_0</ID>952 </input>
<output>
<ID>OUT_0</ID>958 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1053</ID>
<type>AE_DFF_LOW</type>
<position>555.5,-1.5</position>
<input>
<ID>IN_0</ID>1099 </input>
<output>
<ID>OUT_0</ID>1104 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1054</ID>
<type>BA_NAND4</type>
<position>479,117</position>
<input>
<ID>IN_0</ID>1083 </input>
<input>
<ID>IN_1</ID>1082 </input>
<input>
<ID>IN_2</ID>1084 </input>
<input>
<ID>IN_3</ID>1085 </input>
<output>
<ID>OUT</ID>1067 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1055</ID>
<type>AE_SMALL_INVERTER</type>
<position>861,-416</position>
<input>
<ID>IN_0</ID>953 </input>
<output>
<ID>OUT_0</ID>959 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1056</ID>
<type>AE_DFF_LOW</type>
<position>572.5,-1.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1057</ID>
<type>AE_DFF_LOW</type>
<position>588.5,-1.5</position>
<input>
<ID>IN_0</ID>1100 </input>
<output>
<ID>OUT_0</ID>1106 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1058</ID>
<type>AE_SMALL_INVERTER</type>
<position>876,-416</position>
<input>
<ID>IN_0</ID>954 </input>
<output>
<ID>OUT_0</ID>960 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1059</ID>
<type>AE_DFF_LOW</type>
<position>606.5,-1.5</position>
<input>
<ID>IN_0</ID>1101 </input>
<output>
<ID>OUT_0</ID>1107 </output>
<input>
<ID>clear</ID>1062 </input>
<input>
<ID>clock</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1060</ID>
<type>AE_SMALL_INVERTER</type>
<position>891,-416</position>
<input>
<ID>IN_0</ID>955 </input>
<output>
<ID>OUT_0</ID>961 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1061</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>626.5,-11</position>
<input>
<ID>IN_0</ID>1102 </input>
<input>
<ID>IN_1</ID>1103 </input>
<input>
<ID>IN_2</ID>1104 </input>
<input>
<ID>IN_3</ID>1105 </input>
<input>
<ID>IN_4</ID>1106 </input>
<input>
<ID>IN_5</ID>1107 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1062</ID>
<type>AE_SMALL_INVERTER</type>
<position>902.5,-415.5</position>
<input>
<ID>IN_0</ID>956 </input>
<output>
<ID>OUT_0</ID>962 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1063</ID>
<type>AA_INVERTER</type>
<position>514,91.5</position>
<input>
<ID>IN_0</ID>1066 </input>
<output>
<ID>OUT_0</ID>1109 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1064</ID>
<type>AE_SMALL_INVERTER</type>
<position>915.5,-416</position>
<input>
<ID>IN_0</ID>957 </input>
<output>
<ID>OUT_0</ID>963 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1065</ID>
<type>AE_DFF_LOW</type>
<position>396,71.5</position>
<input>
<ID>IN_0</ID>1079 </input>
<output>
<ID>OUT_0</ID>1086 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1066</ID>
<type>AE_SMALL_INVERTER</type>
<position>928.5,-415.5</position>
<input>
<ID>IN_0</ID>958 </input>
<output>
<ID>OUT_0</ID>964 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1067</ID>
<type>AE_DFF_LOW</type>
<position>412.5,71.5</position>
<input>
<ID>IN_0</ID>1081 </input>
<output>
<ID>OUT_0</ID>1087 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1068</ID>
<type>AE_DFF_LOW</type>
<position>427,71.5</position>
<input>
<ID>IN_0</ID>1083 </input>
<output>
<ID>OUT_0</ID>1088 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1069</ID>
<type>AE_DFF_LOW</type>
<position>444,71.5</position>
<input>
<ID>IN_0</ID>1082 </input>
<output>
<ID>OUT_0</ID>1089 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1070</ID>
<type>AE_DFF_LOW</type>
<position>460,71.5</position>
<input>
<ID>IN_0</ID>1084 </input>
<output>
<ID>OUT_0</ID>1090 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1071</ID>
<type>AE_DFF_LOW</type>
<position>478,71.5</position>
<input>
<ID>IN_0</ID>1085 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<input>
<ID>clear</ID>1066 </input>
<input>
<ID>clock</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1072</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>498,62</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1087 </input>
<input>
<ID>IN_2</ID>1088 </input>
<input>
<ID>IN_3</ID>1089 </input>
<input>
<ID>IN_4</ID>1090 </input>
<input>
<ID>IN_5</ID>1091 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1073</ID>
<type>AA_AND2</type>
<position>360.5,102.5</position>
<input>
<ID>IN_0</ID>989 </input>
<input>
<ID>IN_1</ID>996 </input>
<output>
<ID>OUT</ID>1108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1074</ID>
<type>AE_DFF_LOW</type>
<position>304.5,-64.5</position>
<input>
<ID>IN_0</ID>991 </input>
<output>
<ID>OUTINV_0</ID>997 </output>
<output>
<ID>OUT_0</ID>995 </output>
<input>
<ID>clock</ID>993 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1075</ID>
<type>AA_TOGGLE</type>
<position>292,-62.5</position>
<output>
<ID>OUT_0</ID>991 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1076</ID>
<type>AI_XOR2</type>
<position>849,-284.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<input>
<ID>IN_1</ID>1113 </input>
<output>
<ID>OUT</ID>968 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1077</ID>
<type>AI_XOR2</type>
<position>862.5,-284.5</position>
<input>
<ID>IN_0</ID>1103 </input>
<input>
<ID>IN_1</ID>1115 </input>
<output>
<ID>OUT</ID>969 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1078</ID>
<type>AA_AND2</type>
<position>321,-53.5</position>
<input>
<ID>IN_0</ID>995 </input>
<input>
<ID>IN_1</ID>994 </input>
<output>
<ID>OUT</ID>996 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1079</ID>
<type>AI_XOR2</type>
<position>875.5,-284.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>970 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1080</ID>
<type>AA_LABEL</type>
<position>288,-53</position>
<gparam>LABEL_TEXT On/Off Switch</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1081</ID>
<type>AI_XOR2</type>
<position>888.5,-284.5</position>
<input>
<ID>IN_0</ID>1105 </input>
<input>
<ID>IN_1</ID>1119 </input>
<output>
<ID>OUT</ID>971 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1082</ID>
<type>AI_XOR2</type>
<position>901,-285</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1121 </input>
<output>
<ID>OUT</ID>972 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1083</ID>
<type>AE_SMALL_INVERTER</type>
<position>315,-65.5</position>
<input>
<ID>IN_0</ID>997 </input>
<output>
<ID>OUT_0</ID>998 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1084</ID>
<type>AI_XOR2</type>
<position>913.5,-285</position>
<input>
<ID>IN_0</ID>1107 </input>
<input>
<ID>IN_1</ID>1123 </input>
<output>
<ID>OUT</ID>973 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1085</ID>
<type>AA_LABEL</type>
<position>443,-75</position>
<gparam>LABEL_TEXT Default Power</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1086</ID>
<type>AE_DFF_LOW</type>
<position>354.5,-66.5</position>
<input>
<ID>IN_0</ID>992 </input>
<output>
<ID>OUTINV_0</ID>994 </output>
<output>
<ID>OUT_0</ID>1050 </output>
<input>
<ID>clear</ID>998 </input>
<input>
<ID>clock</ID>993 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1087</ID>
<type>BB_CLOCK</type>
<position>339.5,-70</position>
<output>
<ID>CLK</ID>993 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1088</ID>
<type>AA_TOGGLE</type>
<position>735.5,-331</position>
<output>
<ID>OUT_0</ID>1110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1089</ID>
<type>AA_AND2</type>
<position>761.5,-392</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1005 </input>
<output>
<ID>OUT</ID>1124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1090</ID>
<type>AA_AND2</type>
<position>761,-383.5</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1023 </input>
<output>
<ID>OUT</ID>1126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1091</ID>
<type>AA_AND2</type>
<position>760.5,-375</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1024 </input>
<output>
<ID>OUT</ID>1128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1092</ID>
<type>AA_AND2</type>
<position>760,-367</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1093</ID>
<type>AA_AND2</type>
<position>759.5,-358.5</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1026 </input>
<output>
<ID>OUT</ID>1132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1094</ID>
<type>AA_AND2</type>
<position>759.5,-350</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1027 </input>
<output>
<ID>OUT</ID>1134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1095</ID>
<type>AA_LABEL</type>
<position>740.5,-181.5</position>
<gparam>LABEL_TEXT Zone 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1096</ID>
<type>AA_LABEL</type>
<position>743,-318</position>
<gparam>LABEL_TEXT Zone 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1097</ID>
<type>GA_LED</type>
<position>912,-452.5</position>
<input>
<ID>N_in0</ID>1111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1098</ID>
<type>BE_JKFF_LOW_NT</type>
<position>828,-247.5</position>
<input>
<ID>J</ID>1112 </input>
<output>
<ID>Q</ID>1113 </output>
<input>
<ID>clear</ID>1139 </input>
<input>
<ID>clock</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1099</ID>
<type>BE_JKFF_LOW_NT</type>
<position>815,-237.5</position>
<input>
<ID>J</ID>1114 </input>
<output>
<ID>Q</ID>1115 </output>
<input>
<ID>clear</ID>1139 </input>
<input>
<ID>clock</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1100</ID>
<type>BE_JKFF_LOW_NT</type>
<position>802,-226.5</position>
<input>
<ID>J</ID>1116 </input>
<output>
<ID>Q</ID>1117 </output>
<input>
<ID>clear</ID>1139 </input>
<input>
<ID>clock</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1101</ID>
<type>BE_JKFF_LOW_NT</type>
<position>794.5,-217.5</position>
<input>
<ID>J</ID>1118 </input>
<output>
<ID>Q</ID>1119 </output>
<input>
<ID>clear</ID>1139 </input>
<input>
<ID>clock</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1102</ID>
<type>BE_JKFF_LOW_NT</type>
<position>786,-210</position>
<input>
<ID>J</ID>1120 </input>
<output>
<ID>Q</ID>1121 </output>
<input>
<ID>clear</ID>1139 </input>
<input>
<ID>clock</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1103</ID>
<type>BE_JKFF_LOW_NT</type>
<position>777,-202.5</position>
<input>
<ID>J</ID>1122 </input>
<output>
<ID>Q</ID>1123 </output>
<input>
<ID>clear</ID>1139 </input>
<input>
<ID>clock</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1104</ID>
<type>BE_JKFF_LOW_NT</type>
<position>819.5,-394</position>
<input>
<ID>J</ID>1124 </input>
<output>
<ID>Q</ID>1125 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1105</ID>
<type>BE_JKFF_LOW_NT</type>
<position>811.5,-385.5</position>
<input>
<ID>J</ID>1126 </input>
<output>
<ID>Q</ID>1127 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1106</ID>
<type>BE_JKFF_LOW_NT</type>
<position>804.5,-377</position>
<input>
<ID>J</ID>1128 </input>
<output>
<ID>Q</ID>1129 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1107</ID>
<type>BE_JKFF_LOW_NT</type>
<position>795.5,-369</position>
<input>
<ID>J</ID>1130 </input>
<output>
<ID>Q</ID>1131 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1108</ID>
<type>BE_JKFF_LOW_NT</type>
<position>788.5,-360.5</position>
<input>
<ID>J</ID>1132 </input>
<output>
<ID>Q</ID>1133 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1109</ID>
<type>BE_JKFF_LOW_NT</type>
<position>780.5,-352</position>
<input>
<ID>J</ID>1134 </input>
<output>
<ID>Q</ID>1135 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1110</ID>
<type>AA_TOGGLE</type>
<position>810.5,-356</position>
<output>
<ID>OUT_0</ID>1136 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1111</ID>
<type>AA_LABEL</type>
<position>819.5,-353.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1112</ID>
<type>CC_PULSE</type>
<position>773,-344</position>
<output>
<ID>OUT_0</ID>1137 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>1113</ID>
<type>CC_PULSE</type>
<position>769.5,-194.5</position>
<output>
<ID>OUT_0</ID>1138 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>1114</ID>
<type>AA_TOGGLE</type>
<position>835.5,-194.5</position>
<output>
<ID>OUT_0</ID>1139 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1115</ID>
<type>AA_AND4</type>
<position>879,-432.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>961 </input>
<input>
<ID>IN_2</ID>960 </input>
<input>
<ID>IN_3</ID>959 </input>
<output>
<ID>OUT</ID>965 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1116</ID>
<type>AA_AND2</type>
<position>915.5,-431.5</position>
<input>
<ID>IN_0</ID>964 </input>
<input>
<ID>IN_1</ID>963 </input>
<output>
<ID>OUT</ID>966 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1117</ID>
<type>AA_AND2</type>
<position>894.5,-444.5</position>
<input>
<ID>IN_0</ID>966 </input>
<input>
<ID>IN_1</ID>965 </input>
<output>
<ID>OUT</ID>1111 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1118</ID>
<type>AI_XOR2</type>
<position>850,-399.5</position>
<input>
<ID>IN_0</ID>1102 </input>
<input>
<ID>IN_1</ID>1125 </input>
<output>
<ID>OUT</ID>947 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1119</ID>
<type>AI_XOR2</type>
<position>863.5,-399.5</position>
<input>
<ID>IN_0</ID>1103 </input>
<input>
<ID>IN_1</ID>1127 </input>
<output>
<ID>OUT</ID>948 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1120</ID>
<type>AI_XOR2</type>
<position>876.5,-399.5</position>
<input>
<ID>IN_0</ID>1104 </input>
<input>
<ID>IN_1</ID>1129 </input>
<output>
<ID>OUT</ID>949 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1121</ID>
<type>AI_XOR2</type>
<position>889.5,-399.5</position>
<input>
<ID>IN_0</ID>1105 </input>
<input>
<ID>IN_1</ID>1131 </input>
<output>
<ID>OUT</ID>950 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1122</ID>
<type>AI_XOR2</type>
<position>902,-400</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1133 </input>
<output>
<ID>OUT</ID>951 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1123</ID>
<type>AI_XOR2</type>
<position>914.5,-400</position>
<input>
<ID>IN_0</ID>1107 </input>
<input>
<ID>IN_1</ID>1135 </input>
<output>
<ID>OUT</ID>952 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1124</ID>
<type>AE_DFF_LOW</type>
<position>854,-408</position>
<input>
<ID>IN_0</ID>947 </input>
<output>
<ID>OUT_0</ID>953 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1125</ID>
<type>AA_AND2</type>
<position>763,-245.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1005 </input>
<output>
<ID>OUT</ID>1112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1126</ID>
<type>AA_AND2</type>
<position>762.5,-235.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1023 </input>
<output>
<ID>OUT</ID>1114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1127</ID>
<type>AA_AND2</type>
<position>761,-224.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1024 </input>
<output>
<ID>OUT</ID>1116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1128</ID>
<type>AA_AND2</type>
<position>760.5,-215.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1129</ID>
<type>AA_AND2</type>
<position>759.5,-208</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1026 </input>
<output>
<ID>OUT</ID>1120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1130</ID>
<type>AA_AND2</type>
<position>758.5,-200.5</position>
<input>
<ID>IN_0</ID>967 </input>
<input>
<ID>IN_1</ID>1027 </input>
<output>
<ID>OUT</ID>1122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1131</ID>
<type>AA_LABEL</type>
<position>472,-203.5</position>
<gparam>LABEL_TEXT Checking condition for 60</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1132</ID>
<type>AA_TOGGLE</type>
<position>341.5,-64.5</position>
<output>
<ID>OUT_0</ID>992 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1133</ID>
<type>AA_LABEL</type>
<position>673.5,-122.5</position>
<gparam>LABEL_TEXT Problematic Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1134</ID>
<type>BA_NAND4</type>
<position>650.5,-67.5</position>
<input>
<ID>IN_0</ID>1009 </input>
<input>
<ID>IN_1</ID>1013 </input>
<input>
<ID>IN_2</ID>1017 </input>
<input>
<ID>IN_3</ID>1022 </input>
<output>
<ID>OUT</ID>999 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1135</ID>
<type>AE_DFF_LOW</type>
<position>451.5,-137.5</position>
<input>
<ID>IN_0</ID>1000 </input>
<output>
<ID>OUT_0</ID>1005 </output>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1136</ID>
<type>BE_JKFF_LOW_NT</type>
<position>433.5,-93</position>
<input>
<ID>J</ID>1028 </input>
<input>
<ID>K</ID>1030 </input>
<output>
<ID>Q</ID>1000 </output>
<input>
<ID>clear</ID>999 </input>
<input>
<ID>clock</ID>1021 </input>
<output>
<ID>nQ</ID>1001 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1137</ID>
<type>BE_JKFF_LOW_NT</type>
<position>483,-93.5</position>
<input>
<ID>J</ID>1040 </input>
<input>
<ID>K</ID>1041 </input>
<output>
<ID>Q</ID>1004 </output>
<input>
<ID>clear</ID>999 </input>
<input>
<ID>clock</ID>1021 </input>
<output>
<ID>nQ</ID>1007 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1138</ID>
<type>AE_DFF_LOW</type>
<position>494.5,-137</position>
<input>
<ID>IN_0</ID>1004 </input>
<output>
<ID>OUT_0</ID>1023 </output>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1139</ID>
<type>BE_JKFF_LOW_NT</type>
<position>509,-93</position>
<input>
<ID>J</ID>1042 </input>
<input>
<ID>K</ID>1043 </input>
<output>
<ID>Q</ID>1009 </output>
<input>
<ID>clear</ID>999 </input>
<input>
<ID>clock</ID>1021 </input>
<output>
<ID>nQ</ID>1012 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1140</ID>
<type>BE_JKFF_LOW_NT</type>
<position>539,-93.5</position>
<input>
<ID>J</ID>1044 </input>
<input>
<ID>K</ID>1045 </input>
<output>
<ID>Q</ID>1013 </output>
<input>
<ID>clear</ID>999 </input>
<input>
<ID>clock</ID>1021 </input>
<output>
<ID>nQ</ID>1014 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1141</ID>
<type>BE_JKFF_LOW_NT</type>
<position>577.5,-95.5</position>
<input>
<ID>J</ID>1046 </input>
<input>
<ID>K</ID>1047 </input>
<output>
<ID>Q</ID>1017 </output>
<input>
<ID>clear</ID>999 </input>
<input>
<ID>clock</ID>1021 </input>
<output>
<ID>nQ</ID>1018 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1142</ID>
<type>BE_JKFF_LOW_NT</type>
<position>626,-96</position>
<input>
<ID>J</ID>1048 </input>
<input>
<ID>K</ID>1049 </input>
<output>
<ID>Q</ID>1022 </output>
<input>
<ID>clear</ID>999 </input>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1143</ID>
<type>AE_DFF_LOW</type>
<position>524,-137</position>
<input>
<ID>IN_0</ID>1009 </input>
<output>
<ID>OUT_0</ID>1024 </output>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1144</ID>
<type>AA_AND2</type>
<position>450,-84</position>
<input>
<ID>IN_0</ID>1056 </input>
<input>
<ID>IN_1</ID>1000 </input>
<output>
<ID>OUT</ID>1002 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1145</ID>
<type>AE_DFF_LOW</type>
<position>853,-293</position>
<input>
<ID>IN_0</ID>968 </input>
<output>
<ID>OUT_0</ID>974 </output>
<input>
<ID>clock</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1146</ID>
<type>AA_AND2</type>
<position>449,-101.5</position>
<input>
<ID>IN_0</ID>1001 </input>
<input>
<ID>IN_1</ID>1057 </input>
<output>
<ID>OUT</ID>1003 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1147</ID>
<type>AA_AND2</type>
<position>491,-84</position>
<input>
<ID>IN_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1004 </input>
<output>
<ID>OUT</ID>1006 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1148</ID>
<type>AA_AND2</type>
<position>493.5,-102.5</position>
<input>
<ID>IN_0</ID>1007 </input>
<input>
<ID>IN_1</ID>1003 </input>
<output>
<ID>OUT</ID>1008 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1149</ID>
<type>AA_AND2</type>
<position>520.5,-85.5</position>
<input>
<ID>IN_0</ID>1006 </input>
<input>
<ID>IN_1</ID>1009 </input>
<output>
<ID>OUT</ID>1010 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1150</ID>
<type>AA_AND2</type>
<position>523,-104</position>
<input>
<ID>IN_0</ID>1012 </input>
<input>
<ID>IN_1</ID>1008 </input>
<output>
<ID>OUT</ID>1011 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1151</ID>
<type>AA_AND2</type>
<position>547,-86.5</position>
<input>
<ID>IN_0</ID>1010 </input>
<input>
<ID>IN_1</ID>1013 </input>
<output>
<ID>OUT</ID>1015 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1152</ID>
<type>AA_AND2</type>
<position>548.5,-104</position>
<input>
<ID>IN_0</ID>1014 </input>
<input>
<ID>IN_1</ID>1011 </input>
<output>
<ID>OUT</ID>1016 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1153</ID>
<type>AA_AND2</type>
<position>594,-85.5</position>
<input>
<ID>IN_0</ID>1015 </input>
<input>
<ID>IN_1</ID>1017 </input>
<output>
<ID>OUT</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1154</ID>
<type>AA_AND2</type>
<position>594.5,-103</position>
<input>
<ID>IN_0</ID>1018 </input>
<input>
<ID>IN_1</ID>1016 </input>
<output>
<ID>OUT</ID>1020 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1155</ID>
<type>AE_DFF_LOW</type>
<position>552.5,-137</position>
<input>
<ID>IN_0</ID>1013 </input>
<output>
<ID>OUT_0</ID>1025 </output>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1156</ID>
<type>AE_OR2</type>
<position>464,-93.5</position>
<input>
<ID>IN_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1003 </input>
<output>
<ID>OUT</ID>1040 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1157</ID>
<type>AE_DFF_LOW</type>
<position>598.5,-137</position>
<input>
<ID>IN_0</ID>1017 </input>
<output>
<ID>OUT_0</ID>1026 </output>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1158</ID>
<type>AE_OR2</type>
<position>500.5,-92.5</position>
<input>
<ID>IN_0</ID>1006 </input>
<input>
<ID>IN_1</ID>1008 </input>
<output>
<ID>OUT</ID>1043 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1159</ID>
<type>AE_OR2</type>
<position>529,-93</position>
<input>
<ID>IN_0</ID>1010 </input>
<input>
<ID>IN_1</ID>1011 </input>
<output>
<ID>OUT</ID>1044 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1160</ID>
<type>AE_OR2</type>
<position>558,-93.5</position>
<input>
<ID>IN_0</ID>1015 </input>
<input>
<ID>IN_1</ID>1016 </input>
<output>
<ID>OUT</ID>1046 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1161</ID>
<type>AE_OR2</type>
<position>602,-94</position>
<input>
<ID>IN_0</ID>1019 </input>
<input>
<ID>IN_1</ID>1020 </input>
<output>
<ID>OUT</ID>1048 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1162</ID>
<type>AE_DFF_LOW</type>
<position>646.5,-137.5</position>
<input>
<ID>IN_0</ID>1022 </input>
<output>
<ID>OUT_0</ID>1027 </output>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1163</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>650.5,-117</position>
<input>
<ID>IN_0</ID>1000 </input>
<input>
<ID>IN_1</ID>1004 </input>
<input>
<ID>IN_2</ID>1009 </input>
<input>
<ID>IN_3</ID>1013 </input>
<input>
<ID>IN_4</ID>1017 </input>
<input>
<ID>IN_5</ID>1022 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1164</ID>
<type>AE_DFF_LOW</type>
<position>370,-101.5</position>
<input>
<ID>IN_0</ID>1055 </input>
<output>
<ID>OUTINV_0</ID>1057 </output>
<output>
<ID>OUT_0</ID>1056 </output>
<input>
<ID>clear</ID>998 </input>
<input>
<ID>clock</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>947</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>850,-406,850,-402.5</points>
<connection>
<GID>1118</GID>
<name>OUT</name></connection>
<intersection>-406 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>850,-406,851,-406</points>
<connection>
<GID>1124</GID>
<name>IN_0</name></connection>
<intersection>850 0</intersection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>863.5,-406.5,863.5,-402.5</points>
<connection>
<GID>1119</GID>
<name>OUT</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>863.5,-406.5,867,-406.5</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<intersection>863.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>876.5,-406.5,876.5,-402.5</points>
<connection>
<GID>1120</GID>
<name>OUT</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>876.5,-406.5,880.5,-406.5</points>
<connection>
<GID>1039</GID>
<name>IN_0</name></connection>
<intersection>876.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>892.5,-406.5,892.5,-402.5</points>
<intersection>-406.5 1</intersection>
<intersection>-402.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>892.5,-406.5,895.5,-406.5</points>
<connection>
<GID>1044</GID>
<name>IN_0</name></connection>
<intersection>892.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>889.5,-402.5,892.5,-402.5</points>
<connection>
<GID>1121</GID>
<name>OUT</name></connection>
<intersection>892.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>902,-405,902,-403</points>
<connection>
<GID>1122</GID>
<name>OUT</name></connection>
<intersection>-405 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>902,-405,906,-405</points>
<intersection>902 0</intersection>
<intersection>906 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>906,-406.5,906,-405</points>
<connection>
<GID>1050</GID>
<name>IN_0</name></connection>
<intersection>-405 1</intersection></vsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>914.5,-405,914.5,-403</points>
<connection>
<GID>1123</GID>
<name>OUT</name></connection>
<intersection>-405 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>914.5,-405,919,-405</points>
<intersection>914.5 0</intersection>
<intersection>919 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>919,-406.5,919,-405</points>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection>
<intersection>-405 1</intersection></vsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>861,-414,861,-406</points>
<connection>
<GID>1055</GID>
<name>IN_0</name></connection>
<intersection>-406 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>857,-406,861,-406</points>
<connection>
<GID>1124</GID>
<name>OUT_0</name></connection>
<intersection>861 0</intersection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>876,-414,876,-406.5</points>
<connection>
<GID>1058</GID>
<name>IN_0</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>873,-406.5,876,-406.5</points>
<connection>
<GID>1025</GID>
<name>OUT_0</name></connection>
<intersection>876 0</intersection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>891,-414,891,-406.5</points>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>886.5,-406.5,891,-406.5</points>
<connection>
<GID>1039</GID>
<name>OUT_0</name></connection>
<intersection>891 0</intersection></hsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>902.5,-413.5,902.5,-406.5</points>
<connection>
<GID>1062</GID>
<name>IN_0</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>901.5,-406.5,902.5,-406.5</points>
<connection>
<GID>1044</GID>
<name>OUT_0</name></connection>
<intersection>902.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>915.5,-414,915.5,-406.5</points>
<connection>
<GID>1064</GID>
<name>IN_0</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>912,-406.5,915.5,-406.5</points>
<connection>
<GID>1050</GID>
<name>OUT_0</name></connection>
<intersection>915.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>928.5,-413.5,928.5,-406.5</points>
<connection>
<GID>1066</GID>
<name>IN_0</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>925,-406.5,928.5,-406.5</points>
<connection>
<GID>1052</GID>
<name>OUT_0</name></connection>
<intersection>928.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>861,-423.5,861,-418</points>
<connection>
<GID>1055</GID>
<name>OUT_0</name></connection>
<intersection>-423.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>876,-429.5,876,-423.5</points>
<connection>
<GID>1115</GID>
<name>IN_3</name></connection>
<intersection>-423.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>861,-423.5,876,-423.5</points>
<intersection>861 0</intersection>
<intersection>876 1</intersection></hsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>876,-423,876,-418</points>
<connection>
<GID>1058</GID>
<name>OUT_0</name></connection>
<intersection>-423 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>878,-429.5,878,-423</points>
<connection>
<GID>1115</GID>
<name>IN_2</name></connection>
<intersection>-423 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>876,-423,878,-423</points>
<intersection>876 0</intersection>
<intersection>878 1</intersection></hsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>891,-423.5,891,-418</points>
<connection>
<GID>1060</GID>
<name>OUT_0</name></connection>
<intersection>-423.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>880,-429.5,880,-423.5</points>
<connection>
<GID>1115</GID>
<name>IN_1</name></connection>
<intersection>-423.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>880,-423.5,891,-423.5</points>
<intersection>880 1</intersection>
<intersection>891 0</intersection></hsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>902.5,-424.5,902.5,-417.5</points>
<connection>
<GID>1062</GID>
<name>OUT_0</name></connection>
<intersection>-424.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>882,-429.5,882,-424.5</points>
<connection>
<GID>1115</GID>
<name>IN_0</name></connection>
<intersection>-424.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>882,-424.5,902.5,-424.5</points>
<intersection>882 1</intersection>
<intersection>902.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>915.5,-423,915.5,-418</points>
<connection>
<GID>1064</GID>
<name>OUT_0</name></connection>
<intersection>-423 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>914.5,-428.5,914.5,-423</points>
<connection>
<GID>1116</GID>
<name>IN_1</name></connection>
<intersection>-423 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>914.5,-423,915.5,-423</points>
<intersection>914.5 1</intersection>
<intersection>915.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>928.5,-423,928.5,-417.5</points>
<connection>
<GID>1066</GID>
<name>OUT_0</name></connection>
<intersection>-423 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>916.5,-428.5,916.5,-423</points>
<connection>
<GID>1116</GID>
<name>IN_0</name></connection>
<intersection>-423 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>916.5,-423,928.5,-423</points>
<intersection>916.5 1</intersection>
<intersection>928.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>965</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>879,-438.5,879,-435.5</points>
<connection>
<GID>1115</GID>
<name>OUT</name></connection>
<intersection>-438.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>893.5,-441.5,893.5,-438.5</points>
<connection>
<GID>1117</GID>
<name>IN_1</name></connection>
<intersection>-438.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>879,-438.5,893.5,-438.5</points>
<intersection>879 0</intersection>
<intersection>893.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>915.5,-438,915.5,-434.5</points>
<connection>
<GID>1116</GID>
<name>OUT</name></connection>
<intersection>-438 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>895.5,-441.5,895.5,-438</points>
<connection>
<GID>1117</GID>
<name>IN_0</name></connection>
<intersection>-438 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>895.5,-438,915.5,-438</points>
<intersection>895.5 1</intersection>
<intersection>915.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>729,-244.5,729,-187</points>
<connection>
<GID>1013</GID>
<name>OUT_0</name></connection>
<intersection>-244.5 1</intersection>
<intersection>-234.5 3</intersection>
<intersection>-223.5 5</intersection>
<intersection>-214.5 7</intersection>
<intersection>-207 9</intersection>
<intersection>-199.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>729,-244.5,760,-244.5</points>
<connection>
<GID>1125</GID>
<name>IN_0</name></connection>
<intersection>729 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>729,-234.5,759.5,-234.5</points>
<connection>
<GID>1126</GID>
<name>IN_0</name></connection>
<intersection>729 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>729,-223.5,758,-223.5</points>
<connection>
<GID>1127</GID>
<name>IN_0</name></connection>
<intersection>729 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>729,-214.5,757.5,-214.5</points>
<connection>
<GID>1128</GID>
<name>IN_0</name></connection>
<intersection>729 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>729,-207,756.5,-207</points>
<connection>
<GID>1129</GID>
<name>IN_0</name></connection>
<intersection>729 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>729,-199.5,755.5,-199.5</points>
<connection>
<GID>1130</GID>
<name>IN_0</name></connection>
<intersection>729 0</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>849,-291,849,-287.5</points>
<connection>
<GID>1076</GID>
<name>OUT</name></connection>
<intersection>-291 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>849,-291,850,-291</points>
<connection>
<GID>1145</GID>
<name>IN_0</name></connection>
<intersection>849 0</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>862.5,-291.5,862.5,-287.5</points>
<connection>
<GID>1077</GID>
<name>OUT</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>862.5,-291.5,866,-291.5</points>
<connection>
<GID>955</GID>
<name>IN_0</name></connection>
<intersection>862.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>875.5,-291.5,875.5,-287.5</points>
<connection>
<GID>1079</GID>
<name>OUT</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>875.5,-291.5,879.5,-291.5</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<intersection>875.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>891.5,-291.5,891.5,-287.5</points>
<intersection>-291.5 1</intersection>
<intersection>-287.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>891.5,-291.5,894.5,-291.5</points>
<connection>
<GID>971</GID>
<name>IN_0</name></connection>
<intersection>891.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>888.5,-287.5,891.5,-287.5</points>
<connection>
<GID>1081</GID>
<name>OUT</name></connection>
<intersection>891.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>901,-290,901,-288</points>
<connection>
<GID>1082</GID>
<name>OUT</name></connection>
<intersection>-290 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>901,-290,905,-290</points>
<intersection>901 0</intersection>
<intersection>905 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>905,-291.5,905,-290</points>
<connection>
<GID>976</GID>
<name>IN_0</name></connection>
<intersection>-290 1</intersection></vsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>913.5,-290,913.5,-288</points>
<connection>
<GID>1084</GID>
<name>OUT</name></connection>
<intersection>-290 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>913.5,-290,918,-290</points>
<intersection>913.5 0</intersection>
<intersection>918 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>918,-291.5,918,-290</points>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<intersection>-290 1</intersection></vsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>860,-299,860,-291</points>
<connection>
<GID>986</GID>
<name>IN_0</name></connection>
<intersection>-291 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>856,-291,860,-291</points>
<connection>
<GID>1145</GID>
<name>OUT_0</name></connection>
<intersection>860 0</intersection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>875,-299,875,-291.5</points>
<connection>
<GID>989</GID>
<name>IN_0</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>872,-291.5,875,-291.5</points>
<connection>
<GID>955</GID>
<name>OUT_0</name></connection>
<intersection>875 0</intersection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>890,-299,890,-291.5</points>
<connection>
<GID>992</GID>
<name>IN_0</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>885.5,-291.5,890,-291.5</points>
<connection>
<GID>964</GID>
<name>OUT_0</name></connection>
<intersection>890 0</intersection></hsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>901.5,-298.5,901.5,-291.5</points>
<connection>
<GID>994</GID>
<name>IN_0</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>900.5,-291.5,901.5,-291.5</points>
<connection>
<GID>971</GID>
<name>OUT_0</name></connection>
<intersection>901.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>914.5,-299,914.5,-291.5</points>
<connection>
<GID>996</GID>
<name>IN_0</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>911,-291.5,914.5,-291.5</points>
<connection>
<GID>976</GID>
<name>OUT_0</name></connection>
<intersection>914.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>927.5,-298.5,927.5,-291.5</points>
<connection>
<GID>999</GID>
<name>IN_0</name></connection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>924,-291.5,927.5,-291.5</points>
<connection>
<GID>982</GID>
<name>OUT_0</name></connection>
<intersection>927.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>860,-308.5,860,-303</points>
<connection>
<GID>986</GID>
<name>OUT_0</name></connection>
<intersection>-308.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>875,-314.5,875,-308.5</points>
<connection>
<GID>1016</GID>
<name>IN_3</name></connection>
<intersection>-308.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>860,-308.5,875,-308.5</points>
<intersection>860 0</intersection>
<intersection>875 1</intersection></hsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>875,-308,875,-303</points>
<connection>
<GID>989</GID>
<name>OUT_0</name></connection>
<intersection>-308 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>877,-314.5,877,-308</points>
<connection>
<GID>1016</GID>
<name>IN_2</name></connection>
<intersection>-308 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>875,-308,877,-308</points>
<intersection>875 0</intersection>
<intersection>877 1</intersection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>890,-308.5,890,-303</points>
<connection>
<GID>992</GID>
<name>OUT_0</name></connection>
<intersection>-308.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>879,-314.5,879,-308.5</points>
<connection>
<GID>1016</GID>
<name>IN_1</name></connection>
<intersection>-308.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>879,-308.5,890,-308.5</points>
<intersection>879 1</intersection>
<intersection>890 0</intersection></hsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>901.5,-309.5,901.5,-302.5</points>
<connection>
<GID>994</GID>
<name>OUT_0</name></connection>
<intersection>-309.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>881,-314.5,881,-309.5</points>
<connection>
<GID>1016</GID>
<name>IN_0</name></connection>
<intersection>-309.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>881,-309.5,901.5,-309.5</points>
<intersection>881 1</intersection>
<intersection>901.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>914.5,-308,914.5,-303</points>
<connection>
<GID>996</GID>
<name>OUT_0</name></connection>
<intersection>-308 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>913.5,-313.5,913.5,-308</points>
<connection>
<GID>1028</GID>
<name>IN_1</name></connection>
<intersection>-308 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>913.5,-308,914.5,-308</points>
<intersection>913.5 1</intersection>
<intersection>914.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>927.5,-308,927.5,-302.5</points>
<connection>
<GID>999</GID>
<name>OUT_0</name></connection>
<intersection>-308 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>915.5,-313.5,915.5,-308</points>
<connection>
<GID>1028</GID>
<name>IN_0</name></connection>
<intersection>-308 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>915.5,-308,927.5,-308</points>
<intersection>915.5 1</intersection>
<intersection>927.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>878,-323.5,878,-320.5</points>
<connection>
<GID>1016</GID>
<name>OUT</name></connection>
<intersection>-323.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>892.5,-326.5,892.5,-323.5</points>
<connection>
<GID>1031</GID>
<name>IN_1</name></connection>
<intersection>-323.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>878,-323.5,892.5,-323.5</points>
<intersection>878 0</intersection>
<intersection>892.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>914.5,-323,914.5,-319.5</points>
<connection>
<GID>1028</GID>
<name>OUT</name></connection>
<intersection>-323 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>894.5,-326.5,894.5,-323</points>
<connection>
<GID>1031</GID>
<name>IN_0</name></connection>
<intersection>-323 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>894.5,-323,914.5,-323</points>
<intersection>894.5 1</intersection>
<intersection>914.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,122,368,126.5</points>
<connection>
<GID>1038</GID>
<name>IN_1</name></connection>
<intersection>126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358.5,126.5,368,126.5</points>
<connection>
<GID>1020</GID>
<name>OUT_0</name></connection>
<intersection>368 0</intersection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,103.5,356.5,116</points>
<intersection>103.5 1</intersection>
<intersection>116 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356.5,103.5,357.5,103.5</points>
<connection>
<GID>1073</GID>
<name>IN_0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,116,369,116</points>
<connection>
<GID>1038</GID>
<name>OUT</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>946,-332.5,946,131</points>
<intersection>-332.5 4</intersection>
<intersection>131 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>370,131,946,131</points>
<intersection>370 5</intersection>
<intersection>946 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>893.5,-332.5,946,-332.5</points>
<connection>
<GID>1031</GID>
<name>OUT</name></connection>
<intersection>946 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>370,122,370,131</points>
<connection>
<GID>1038</GID>
<name>IN_0</name></connection>
<intersection>131 3</intersection></vsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>294,-62.5,301.5,-62.5</points>
<connection>
<GID>1075</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1074</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343.5,-64.5,351.5,-64.5</points>
<connection>
<GID>1132</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1086</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347.5,-73,347.5,-67.5</points>
<intersection>-73 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347.5,-67.5,351.5,-67.5</points>
<connection>
<GID>1086</GID>
<name>clock</name></connection>
<intersection>347.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-73,347.5,-73</points>
<intersection>301.5 3</intersection>
<intersection>343.5 4</intersection>
<intersection>347.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>301.5,-73,301.5,-65.5</points>
<connection>
<GID>1074</GID>
<name>clock</name></connection>
<intersection>-73 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>343.5,-73,343.5,-70</points>
<connection>
<GID>1087</GID>
<name>CLK</name></connection>
<intersection>-73 2</intersection></vsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,-76.5,322,-56.5</points>
<connection>
<GID>1078</GID>
<name>IN_1</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-76.5,357.5,-76.5</points>
<intersection>322 0</intersection>
<intersection>357.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>357.5,-76.5,357.5,-67.5</points>
<connection>
<GID>1086</GID>
<name>OUTINV_0</name></connection>
<intersection>-76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-62.5,320,-56.5</points>
<connection>
<GID>1078</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>307.5,-62.5,320,-62.5</points>
<connection>
<GID>1074</GID>
<name>OUT_0</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-50.5,321,101.5</points>
<connection>
<GID>1078</GID>
<name>OUT</name></connection>
<intersection>101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,101.5,357.5,101.5</points>
<connection>
<GID>1073</GID>
<name>IN_1</name></connection>
<intersection>321 0</intersection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307.5,-65.5,313,-65.5</points>
<connection>
<GID>1074</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>1083</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-105.5,354.5,-70.5</points>
<connection>
<GID>1086</GID>
<name>clear</name></connection>
<intersection>-105.5 3</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-78,354.5,-78</points>
<intersection>317 2</intersection>
<intersection>354.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>317,-78,317,-65.5</points>
<connection>
<GID>1083</GID>
<name>OUT_0</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>354.5,-105.5,370,-105.5</points>
<connection>
<GID>1164</GID>
<name>clear</name></connection>
<intersection>354.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>658.5,-123,658.5,-67.5</points>
<intersection>-123 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653.5,-67.5,658.5,-67.5</points>
<connection>
<GID>1134</GID>
<name>OUT</name></connection>
<intersection>658.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>433.5,-123,658.5,-123</points>
<intersection>433.5 15</intersection>
<intersection>483 14</intersection>
<intersection>509 10</intersection>
<intersection>539 18</intersection>
<intersection>577.5 16</intersection>
<intersection>626 17</intersection>
<intersection>658.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>509,-123,509,-97</points>
<connection>
<GID>1139</GID>
<name>clear</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>483,-123,483,-97.5</points>
<connection>
<GID>1137</GID>
<name>clear</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>433.5,-123,433.5,-97</points>
<connection>
<GID>1136</GID>
<name>clear</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>577.5,-123,577.5,-99.5</points>
<connection>
<GID>1141</GID>
<name>clear</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>626,-123,626,-100</points>
<connection>
<GID>1142</GID>
<name>clear</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>539,-123,539,-97.5</points>
<connection>
<GID>1140</GID>
<name>clear</name></connection>
<intersection>-123 2</intersection></vsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442.5,-135.5,442.5,-85</points>
<intersection>-135.5 8</intersection>
<intersection>-129.5 5</intersection>
<intersection>-120 3</intersection>
<intersection>-91 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,-85,447,-85</points>
<connection>
<GID>1144</GID>
<name>IN_1</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436.5,-91,442.5,-91</points>
<connection>
<GID>1136</GID>
<name>Q</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>442.5,-120,645.5,-120</points>
<connection>
<GID>1163</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>442.5,-129.5,461.5,-129.5</points>
<intersection>442.5 0</intersection>
<intersection>461.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>461.5,-162,461.5,-129.5</points>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<intersection>-129.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>442.5,-135.5,448.5,-135.5</points>
<connection>
<GID>1135</GID>
<name>IN_0</name></connection>
<intersection>442.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1001</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438.5,-100.5,438.5,-95</points>
<intersection>-100.5 3</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>436.5,-95,438.5,-95</points>
<connection>
<GID>1136</GID>
<name>nQ</name></connection>
<intersection>438.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>438.5,-100.5,446,-100.5</points>
<connection>
<GID>1146</GID>
<name>IN_0</name></connection>
<intersection>438.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-92.5,457,-83</points>
<intersection>-92.5 1</intersection>
<intersection>-84 2</intersection>
<intersection>-83 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>457,-92.5,461,-92.5</points>
<connection>
<GID>1156</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>453,-84,457,-84</points>
<connection>
<GID>1144</GID>
<name>OUT</name></connection>
<intersection>457 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>457,-83,488,-83</points>
<connection>
<GID>1147</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment></shape></wire>
<wire>
<ID>1003</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,-103.5,457.5,-94.5</points>
<intersection>-103.5 2</intersection>
<intersection>-101.5 3</intersection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>457.5,-94.5,461,-94.5</points>
<connection>
<GID>1156</GID>
<name>IN_1</name></connection>
<intersection>457.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>457.5,-103.5,490.5,-103.5</points>
<connection>
<GID>1148</GID>
<name>IN_1</name></connection>
<intersection>457.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>452,-101.5,457.5,-101.5</points>
<connection>
<GID>1146</GID>
<name>OUT</name></connection>
<intersection>457.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>487,-161.5,487,-85</points>
<intersection>-161.5 9</intersection>
<intersection>-135 5</intersection>
<intersection>-119 3</intersection>
<intersection>-91.5 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-85,488,-85</points>
<connection>
<GID>1147</GID>
<name>IN_1</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>486,-91.5,487,-91.5</points>
<connection>
<GID>1137</GID>
<name>Q</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>487,-119,645.5,-119</points>
<connection>
<GID>1163</GID>
<name>IN_1</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>487,-135,491.5,-135</points>
<connection>
<GID>1138</GID>
<name>IN_0</name></connection>
<intersection>487 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>474,-161.5,487,-161.5</points>
<intersection>474 10</intersection>
<intersection>487 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>474,-163,474,-161.5</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<intersection>-161.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457.5,-393,457.5,-135.5</points>
<intersection>-393 12</intersection>
<intersection>-247 5</intersection>
<intersection>-150.5 10</intersection>
<intersection>-135.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454.5,-135.5,457.5,-135.5</points>
<connection>
<GID>1135</GID>
<name>OUT_0</name></connection>
<intersection>457.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>457.5,-247,760,-247</points>
<intersection>457.5 0</intersection>
<intersection>760 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>760,-247,760,-246.5</points>
<connection>
<GID>1125</GID>
<name>IN_1</name></connection>
<intersection>-247 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>457.5,-150.5,665,-150.5</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<intersection>457.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>457.5,-393,758.5,-393</points>
<connection>
<GID>1089</GID>
<name>IN_1</name></connection>
<intersection>457.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495.5,-84.5,495.5,-84</points>
<intersection>-84.5 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>494,-84,495.5,-84</points>
<connection>
<GID>1147</GID>
<name>OUT</name></connection>
<intersection>495.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495.5,-84.5,517.5,-84.5</points>
<connection>
<GID>1149</GID>
<name>IN_0</name></connection>
<intersection>495.5 0</intersection>
<intersection>497.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>497.5,-91.5,497.5,-84.5</points>
<connection>
<GID>1158</GID>
<name>IN_0</name></connection>
<intersection>-84.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488.5,-101.5,488.5,-95.5</points>
<intersection>-101.5 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>486,-95.5,488.5,-95.5</points>
<connection>
<GID>1137</GID>
<name>nQ</name></connection>
<intersection>488.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>488.5,-101.5,490.5,-101.5</points>
<connection>
<GID>1148</GID>
<name>IN_0</name></connection>
<intersection>488.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-105,497,-93.5</points>
<intersection>-105 3</intersection>
<intersection>-102.5 1</intersection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>496.5,-102.5,497,-102.5</points>
<connection>
<GID>1148</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-93.5,497.5,-93.5</points>
<connection>
<GID>1158</GID>
<name>IN_1</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>497,-105,520,-105</points>
<connection>
<GID>1150</GID>
<name>IN_1</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-162,514,-64.5</points>
<intersection>-162 13</intersection>
<intersection>-135 9</intersection>
<intersection>-118 2</intersection>
<intersection>-91 1</intersection>
<intersection>-86.5 5</intersection>
<intersection>-64.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-91,514,-91</points>
<connection>
<GID>1139</GID>
<name>Q</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,-118,645.5,-118</points>
<connection>
<GID>1163</GID>
<name>IN_2</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>514,-86.5,517.5,-86.5</points>
<connection>
<GID>1149</GID>
<name>IN_1</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>514,-64.5,647.5,-64.5</points>
<connection>
<GID>1134</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>514,-135,521,-135</points>
<connection>
<GID>1143</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>514,-162,538,-162</points>
<connection>
<GID>974</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>523.5,-85.5,544,-85.5</points>
<connection>
<GID>1149</GID>
<name>OUT</name></connection>
<connection>
<GID>1151</GID>
<name>IN_0</name></connection>
<intersection>526 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>526,-92,526,-85.5</points>
<connection>
<GID>1159</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>526,-105,526,-94</points>
<connection>
<GID>1159</GID>
<name>IN_1</name></connection>
<connection>
<GID>1150</GID>
<name>OUT</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>526,-105,545.5,-105</points>
<connection>
<GID>1152</GID>
<name>IN_1</name></connection>
<intersection>526 0</intersection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515.5,-103,515.5,-95</points>
<intersection>-103 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512,-95,515.5,-95</points>
<connection>
<GID>1139</GID>
<name>nQ</name></connection>
<intersection>515.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515.5,-103,520,-103</points>
<connection>
<GID>1150</GID>
<name>IN_0</name></connection>
<intersection>515.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542,-135,542,-66.5</points>
<connection>
<GID>1140</GID>
<name>Q</name></connection>
<intersection>-135 10</intersection>
<intersection>-117 2</intersection>
<intersection>-87.5 6</intersection>
<intersection>-66.5 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>542,-117,645.5,-117</points>
<connection>
<GID>1163</GID>
<name>IN_3</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>542,-87.5,544,-87.5</points>
<connection>
<GID>1151</GID>
<name>IN_1</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>542,-66.5,647.5,-66.5</points>
<connection>
<GID>1134</GID>
<name>IN_1</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>542,-135,549.5,-135</points>
<connection>
<GID>1155</GID>
<name>IN_0</name></connection>
<intersection>542 0</intersection>
<intersection>545 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>545,-162,545,-135</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<intersection>-135 10</intersection></vsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543,-103,543,-95.5</points>
<intersection>-103 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>542,-95.5,543,-95.5</points>
<connection>
<GID>1140</GID>
<name>nQ</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>543,-103,545.5,-103</points>
<connection>
<GID>1152</GID>
<name>IN_0</name></connection>
<intersection>543 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>553,-92.5,553,-84.5</points>
<intersection>-92.5 2</intersection>
<intersection>-86.5 1</intersection>
<intersection>-84.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>550,-86.5,553,-86.5</points>
<connection>
<GID>1151</GID>
<name>OUT</name></connection>
<intersection>553 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553,-92.5,555,-92.5</points>
<connection>
<GID>1160</GID>
<name>IN_0</name></connection>
<intersection>553 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>553,-84.5,591,-84.5</points>
<connection>
<GID>1153</GID>
<name>IN_0</name></connection>
<intersection>553 0</intersection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>553.5,-104,553.5,-94.5</points>
<intersection>-104 1</intersection>
<intersection>-94.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>551.5,-104,591.5,-104</points>
<connection>
<GID>1152</GID>
<name>OUT</name></connection>
<connection>
<GID>1154</GID>
<name>IN_1</name></connection>
<intersection>553.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>553.5,-94.5,555,-94.5</points>
<connection>
<GID>1160</GID>
<name>IN_1</name></connection>
<intersection>553.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-161.5,585.5,-68.5</points>
<intersection>-161.5 14</intersection>
<intersection>-135 9</intersection>
<intersection>-116 3</intersection>
<intersection>-93.5 1</intersection>
<intersection>-86.5 10</intersection>
<intersection>-68.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>580.5,-93.5,585.5,-93.5</points>
<connection>
<GID>1141</GID>
<name>Q</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>585.5,-116,645.5,-116</points>
<connection>
<GID>1163</GID>
<name>IN_4</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>585.5,-68.5,647.5,-68.5</points>
<connection>
<GID>1134</GID>
<name>IN_2</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>585.5,-135,595.5,-135</points>
<connection>
<GID>1157</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>585.5,-86.5,591,-86.5</points>
<connection>
<GID>1153</GID>
<name>IN_1</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>585.5,-161.5,602.5,-161.5</points>
<connection>
<GID>977</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583,-102,583,-97.5</points>
<intersection>-102 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>580.5,-97.5,583,-97.5</points>
<connection>
<GID>1141</GID>
<name>nQ</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583,-102,591.5,-102</points>
<connection>
<GID>1154</GID>
<name>IN_0</name></connection>
<intersection>583 0</intersection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>598,-93,598,-85.5</points>
<intersection>-93 2</intersection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597,-85.5,598,-85.5</points>
<connection>
<GID>1153</GID>
<name>OUT</name></connection>
<intersection>598 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>598,-93,599,-93</points>
<connection>
<GID>1161</GID>
<name>IN_0</name></connection>
<intersection>598 0</intersection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>598,-103,598,-95</points>
<intersection>-103 1</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597.5,-103,598,-103</points>
<connection>
<GID>1154</GID>
<name>OUT</name></connection>
<intersection>598 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>598,-95,599,-95</points>
<connection>
<GID>1161</GID>
<name>IN_1</name></connection>
<intersection>598 0</intersection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>405,-112.5,623,-112.5</points>
<intersection>405 16</intersection>
<intersection>422.5 13</intersection>
<intersection>479.5 12</intersection>
<intersection>505 6</intersection>
<intersection>533 7</intersection>
<intersection>571 11</intersection>
<intersection>623 28</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>505,-112.5,505,-93</points>
<intersection>-112.5 1</intersection>
<intersection>-93 19</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>533,-112.5,533,-93.5</points>
<intersection>-112.5 1</intersection>
<intersection>-93.5 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>571,-112.5,571,-95.5</points>
<intersection>-112.5 1</intersection>
<intersection>-95.5 18</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>479.5,-112.5,479.5,-93.5</points>
<intersection>-112.5 1</intersection>
<intersection>-93.5 22</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>422.5,-112.5,422.5,-93</points>
<intersection>-112.5 1</intersection>
<intersection>-93 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>533,-93.5,536,-93.5</points>
<connection>
<GID>1140</GID>
<name>clock</name></connection>
<intersection>533 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>422.5,-93,430.5,-93</points>
<connection>
<GID>1136</GID>
<name>clock</name></connection>
<intersection>422.5 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>405,-142,405,-112.5</points>
<intersection>-142 17</intersection>
<intersection>-113 37</intersection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>405,-142,643.5,-142</points>
<intersection>405 16</intersection>
<intersection>448.5 34</intersection>
<intersection>491.5 25</intersection>
<intersection>521 26</intersection>
<intersection>549.5 24</intersection>
<intersection>594.5 23</intersection>
<intersection>643.5 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>571,-95.5,574.5,-95.5</points>
<connection>
<GID>1141</GID>
<name>clock</name></connection>
<intersection>571 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>505,-93,506,-93</points>
<connection>
<GID>1139</GID>
<name>clock</name></connection>
<intersection>505 6</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>479.5,-93.5,480,-93.5</points>
<connection>
<GID>1137</GID>
<name>clock</name></connection>
<intersection>479.5 12</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>594.5,-142,594.5,-138</points>
<intersection>-142 17</intersection>
<intersection>-138 36</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>549.5,-142,549.5,-138</points>
<connection>
<GID>1155</GID>
<name>clock</name></connection>
<intersection>-142 17</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>491.5,-142,491.5,-138</points>
<connection>
<GID>1138</GID>
<name>clock</name></connection>
<intersection>-142 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>521,-142,521,-138</points>
<connection>
<GID>1143</GID>
<name>clock</name></connection>
<intersection>-142 17</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>623,-112.5,623,-96</points>
<connection>
<GID>1142</GID>
<name>clock</name></connection>
<intersection>-112.5 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>448.5,-142,448.5,-138.5</points>
<connection>
<GID>1135</GID>
<name>clock</name></connection>
<intersection>-142 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>643.5,-142,643.5,-138.5</points>
<connection>
<GID>1162</GID>
<name>clock</name></connection>
<intersection>-142 17</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>594.5,-138,595.5,-138</points>
<connection>
<GID>1157</GID>
<name>clock</name></connection>
<intersection>594.5 23</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>364,-113,405,-113</points>
<connection>
<GID>954</GID>
<name>OUT</name></connection>
<intersection>366.5 38</intersection>
<intersection>405 16</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>366.5,-113,366.5,-102.5</points>
<intersection>-113 37</intersection>
<intersection>-102.5 39</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>366.5,-102.5,367,-102.5</points>
<connection>
<GID>1164</GID>
<name>clock</name></connection>
<intersection>366.5 38</intersection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638,-161,638,-70.5</points>
<intersection>-161 9</intersection>
<intersection>-135.5 13</intersection>
<intersection>-115 2</intersection>
<intersection>-94 11</intersection>
<intersection>-70.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>638,-115,645.5,-115</points>
<connection>
<GID>1163</GID>
<name>IN_5</name></connection>
<intersection>638 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>638,-70.5,647.5,-70.5</points>
<connection>
<GID>1134</GID>
<name>IN_3</name></connection>
<intersection>638 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>608,-161,638,-161</points>
<connection>
<GID>978</GID>
<name>IN_0</name></connection>
<intersection>638 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>629,-94,638,-94</points>
<connection>
<GID>1142</GID>
<name>Q</name></connection>
<intersection>638 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>638,-135.5,643.5,-135.5</points>
<connection>
<GID>1162</GID>
<name>IN_0</name></connection>
<intersection>638 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>499,-384.5,499,-135</points>
<intersection>-384.5 16</intersection>
<intersection>-236.5 11</intersection>
<intersection>-149.5 14</intersection>
<intersection>-135 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>497.5,-135,499,-135</points>
<connection>
<GID>1138</GID>
<name>OUT_0</name></connection>
<intersection>499 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>499,-236.5,759.5,-236.5</points>
<connection>
<GID>1126</GID>
<name>IN_1</name></connection>
<intersection>499 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>499,-149.5,665,-149.5</points>
<connection>
<GID>951</GID>
<name>IN_1</name></connection>
<intersection>499 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>499,-384.5,758,-384.5</points>
<connection>
<GID>1090</GID>
<name>IN_1</name></connection>
<intersection>499 3</intersection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>528.5,-376,528.5,-135</points>
<intersection>-376 14</intersection>
<intersection>-225.5 7</intersection>
<intersection>-148.5 12</intersection>
<intersection>-135 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>527,-135,528.5,-135</points>
<connection>
<GID>1143</GID>
<name>OUT_0</name></connection>
<intersection>528.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>528.5,-225.5,758,-225.5</points>
<connection>
<GID>1127</GID>
<name>IN_1</name></connection>
<intersection>528.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>528.5,-148.5,665,-148.5</points>
<connection>
<GID>951</GID>
<name>IN_2</name></connection>
<intersection>528.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>528.5,-376,757.5,-376</points>
<connection>
<GID>1091</GID>
<name>IN_1</name></connection>
<intersection>528.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>555.5,-368,555.5,-135</points>
<connection>
<GID>1155</GID>
<name>OUT_0</name></connection>
<intersection>-368 17</intersection>
<intersection>-216.5 7</intersection>
<intersection>-147.5 15</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>555.5,-216.5,757.5,-216.5</points>
<connection>
<GID>1128</GID>
<name>IN_1</name></connection>
<intersection>555.5 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>555.5,-147.5,665,-147.5</points>
<connection>
<GID>951</GID>
<name>IN_3</name></connection>
<intersection>555.5 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>555.5,-368,757,-368</points>
<connection>
<GID>1092</GID>
<name>IN_1</name></connection>
<intersection>555.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>613.5,-359.5,613.5,-135</points>
<intersection>-359.5 12</intersection>
<intersection>-209 5</intersection>
<intersection>-146.5 10</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>601.5,-135,613.5,-135</points>
<connection>
<GID>1157</GID>
<name>OUT_0</name></connection>
<intersection>613.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>613.5,-209,756.5,-209</points>
<connection>
<GID>1129</GID>
<name>IN_1</name></connection>
<intersection>613.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>613.5,-146.5,665,-146.5</points>
<connection>
<GID>951</GID>
<name>IN_4</name></connection>
<intersection>613.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>613.5,-359.5,756.5,-359.5</points>
<connection>
<GID>1093</GID>
<name>IN_1</name></connection>
<intersection>613.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>656.5,-351,656.5,-135.5</points>
<intersection>-351 18</intersection>
<intersection>-201.5 10</intersection>
<intersection>-145.5 16</intersection>
<intersection>-135.5 13</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>656.5,-201.5,755.5,-201.5</points>
<connection>
<GID>1130</GID>
<name>IN_1</name></connection>
<intersection>656.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>649.5,-135.5,656.5,-135.5</points>
<connection>
<GID>1162</GID>
<name>OUT_0</name></connection>
<intersection>656.5 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>656.5,-145.5,665,-145.5</points>
<connection>
<GID>951</GID>
<name>IN_5</name></connection>
<intersection>656.5 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>656.5,-351,756.5,-351</points>
<connection>
<GID>1094</GID>
<name>IN_1</name></connection>
<intersection>656.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-91,427.5,-78.5</points>
<intersection>-91 8</intersection>
<intersection>-78.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>419,-78.5,427.5,-78.5</points>
<intersection>419 9</intersection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>427.5,-91,430.5,-91</points>
<connection>
<GID>1136</GID>
<name>J</name></connection>
<intersection>427.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>419,-79,419,-67</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<intersection>-78.5 6</intersection>
<intersection>-67 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>378,-67,419,-67</points>
<intersection>378 14</intersection>
<intersection>419 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>378,-70.5,378,-67</points>
<intersection>-70.5 15</intersection>
<intersection>-67 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>367.5,-70.5,378,-70.5</points>
<connection>
<GID>980</GID>
<name>OUT</name></connection>
<intersection>378 14</intersection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>412.5,-71.5,610.5,-71.5</points>
<intersection>412.5 7</intersection>
<intersection>468 6</intersection>
<intersection>504.5 10</intersection>
<intersection>533 12</intersection>
<intersection>563 14</intersection>
<intersection>610.5 16</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>468,-76.5,468,-71.5</points>
<connection>
<GID>965</GID>
<name>IN_1</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>412.5,-78.5,412.5,-71.5</points>
<intersection>-78.5 20</intersection>
<intersection>-71.5 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>504.5,-76,504.5,-71.5</points>
<connection>
<GID>966</GID>
<name>IN_1</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>533,-76.5,533,-71.5</points>
<connection>
<GID>967</GID>
<name>IN_1</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>563,-76.5,563,-71.5</points>
<connection>
<GID>968</GID>
<name>IN_1</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>610.5,-74.5,610.5,-71.5</points>
<connection>
<GID>969</GID>
<name>IN_1</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>382,-78.5,417,-78.5</points>
<intersection>382 23</intersection>
<intersection>412.5 7</intersection>
<intersection>417 26</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>382,-214,382,-78.5</points>
<intersection>-214 24</intersection>
<intersection>-78.5 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>382,-214,446,-214</points>
<intersection>382 23</intersection>
<intersection>446 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>446,-214,446,-213</points>
<connection>
<GID>970</GID>
<name>OUT</name></connection>
<intersection>-214 24</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>417,-79,417,-78.5</points>
<connection>
<GID>963</GID>
<name>IN_1</name></connection>
<intersection>-78.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>418,-95,418,-85</points>
<connection>
<GID>963</GID>
<name>OUT</name></connection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>418,-95,430.5,-95</points>
<connection>
<GID>1136</GID>
<name>K</name></connection>
<intersection>418 0</intersection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466.5,-185,466.5,-173.5</points>
<connection>
<GID>957</GID>
<name>IN_1</name></connection>
<intersection>-173.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>461.5,-173.5,461.5,-168</points>
<connection>
<GID>972</GID>
<name>OUT_0</name></connection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>461.5,-173.5,466.5,-173.5</points>
<intersection>461.5 1</intersection>
<intersection>466.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468.5,-185,468.5,-173.5</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<intersection>-173.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>474,-173.5,474,-169</points>
<connection>
<GID>973</GID>
<name>OUT_0</name></connection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>468.5,-173.5,474,-173.5</points>
<intersection>468.5 0</intersection>
<intersection>474 1</intersection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445,-207,445,-194.5</points>
<connection>
<GID>970</GID>
<name>IN_2</name></connection>
<intersection>-194.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>467.5,-194.5,467.5,-191</points>
<connection>
<GID>957</GID>
<name>OUT</name></connection>
<intersection>-194.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>445,-194.5,467.5,-194.5</points>
<intersection>445 0</intersection>
<intersection>467.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542.5,-171.5,542.5,-169.5</points>
<connection>
<GID>960</GID>
<name>IN_0</name></connection>
<intersection>-169.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>545,-169.5,545,-168</points>
<connection>
<GID>975</GID>
<name>OUT_0</name></connection>
<intersection>-169.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>542.5,-169.5,545,-169.5</points>
<intersection>542.5 0</intersection>
<intersection>545 1</intersection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-171.5,540.5,-169.5</points>
<connection>
<GID>960</GID>
<name>IN_1</name></connection>
<intersection>-169.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>538,-169.5,538,-168</points>
<connection>
<GID>974</GID>
<name>OUT_0</name></connection>
<intersection>-169.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>538,-169.5,540.5,-169.5</points>
<intersection>538 1</intersection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>447,-207,447,-196.5</points>
<connection>
<GID>970</GID>
<name>IN_1</name></connection>
<intersection>-196.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>541.5,-196.5,541.5,-177.5</points>
<connection>
<GID>960</GID>
<name>OUT</name></connection>
<intersection>-196.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>447,-196.5,541.5,-196.5</points>
<intersection>447 0</intersection>
<intersection>541.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-170,605.5,-168.5</points>
<connection>
<GID>962</GID>
<name>IN_0</name></connection>
<intersection>-168.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>608,-168.5,608,-167</points>
<connection>
<GID>978</GID>
<name>OUT_0</name></connection>
<intersection>-168.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>605.5,-168.5,608,-168.5</points>
<intersection>605.5 0</intersection>
<intersection>608 1</intersection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603.5,-170,603.5,-168.5</points>
<connection>
<GID>962</GID>
<name>IN_1</name></connection>
<intersection>-168.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>602.5,-168.5,602.5,-167.5</points>
<connection>
<GID>977</GID>
<name>OUT_0</name></connection>
<intersection>-168.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>602.5,-168.5,603.5,-168.5</points>
<intersection>602.5 1</intersection>
<intersection>603.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449,-207,449,-199</points>
<connection>
<GID>970</GID>
<name>IN_0</name></connection>
<intersection>-199 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>604.5,-199,604.5,-176</points>
<connection>
<GID>962</GID>
<name>OUT</name></connection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>449,-199,604.5,-199</points>
<intersection>449 0</intersection>
<intersection>604.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477.5,-93.5,477.5,-76</points>
<intersection>-93.5 2</intersection>
<intersection>-91.5 1</intersection>
<intersection>-76 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477.5,-91.5,480,-91.5</points>
<connection>
<GID>1137</GID>
<name>J</name></connection>
<intersection>477.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>467,-93.5,477.5,-93.5</points>
<connection>
<GID>1156</GID>
<name>OUT</name></connection>
<intersection>477.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>470,-76,477.5,-76</points>
<intersection>470 4</intersection>
<intersection>477.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>470,-76.5,470,-76</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>-76 3</intersection></vsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469,-95.5,469,-82.5</points>
<connection>
<GID>965</GID>
<name>OUT</name></connection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>469,-95.5,480,-95.5</points>
<connection>
<GID>1137</GID>
<name>K</name></connection>
<intersection>469 0</intersection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,-91,505.5,-82</points>
<connection>
<GID>966</GID>
<name>OUT</name></connection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505.5,-91,506,-91</points>
<connection>
<GID>1139</GID>
<name>J</name></connection>
<intersection>505.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,-83.5,513,-76</points>
<intersection>-83.5 1</intersection>
<intersection>-76 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503.5,-83.5,513,-83.5</points>
<intersection>503.5 4</intersection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>506.5,-76,513,-76</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>513 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>503.5,-95,503.5,-83.5</points>
<connection>
<GID>1158</GID>
<name>OUT</name></connection>
<intersection>-95 6</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>503.5,-95,506,-95</points>
<connection>
<GID>1139</GID>
<name>K</name></connection>
<intersection>503.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>532,-84,538.5,-84</points>
<intersection>532 3</intersection>
<intersection>538.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>532,-93,532,-84</points>
<connection>
<GID>1159</GID>
<name>OUT</name></connection>
<intersection>-91.5 7</intersection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>538.5,-84,538.5,-76.5</points>
<intersection>-84 1</intersection>
<intersection>-76.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>535,-76.5,538.5,-76.5</points>
<connection>
<GID>967</GID>
<name>IN_0</name></connection>
<intersection>538.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>532,-91.5,536,-91.5</points>
<connection>
<GID>1140</GID>
<name>J</name></connection>
<intersection>532 3</intersection></hsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534,-95.5,534,-82.5</points>
<connection>
<GID>967</GID>
<name>OUT</name></connection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,-95.5,536,-95.5</points>
<connection>
<GID>1140</GID>
<name>K</name></connection>
<intersection>534 0</intersection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>561,-93.5,574.5,-93.5</points>
<connection>
<GID>1160</GID>
<name>OUT</name></connection>
<connection>
<GID>1141</GID>
<name>J</name></connection>
<intersection>567.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>567.5,-93.5,567.5,-75.5</points>
<intersection>-93.5 1</intersection>
<intersection>-75.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>565,-75.5,567.5,-75.5</points>
<intersection>565 6</intersection>
<intersection>567.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>565,-76.5,565,-75.5</points>
<connection>
<GID>968</GID>
<name>IN_0</name></connection>
<intersection>-75.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564,-97.5,564,-82.5</points>
<connection>
<GID>968</GID>
<name>OUT</name></connection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>564,-97.5,574.5,-97.5</points>
<connection>
<GID>1141</GID>
<name>K</name></connection>
<intersection>564 0</intersection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>605,-94,623,-94</points>
<connection>
<GID>1161</GID>
<name>OUT</name></connection>
<connection>
<GID>1142</GID>
<name>J</name></connection>
<intersection>613 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>613,-94,613,-73</points>
<intersection>-94 1</intersection>
<intersection>-73 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>612.5,-73,613,-73</points>
<intersection>612.5 15</intersection>
<intersection>613 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>612.5,-74.5,612.5,-73</points>
<connection>
<GID>969</GID>
<name>IN_0</name></connection>
<intersection>-73 8</intersection></vsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>611.5,-98,611.5,-80.5</points>
<connection>
<GID>969</GID>
<name>OUT</name></connection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>611.5,-98,623,-98</points>
<connection>
<GID>1142</GID>
<name>K</name></connection>
<intersection>611.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>357.5,-64.5,366.5,-64.5</points>
<connection>
<GID>980</GID>
<name>IN_1</name></connection>
<connection>
<GID>1086</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368.5,-64.5,368.5,-63.5</points>
<connection>
<GID>980</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>374.5,-63.5,374.5,-62</points>
<connection>
<GID>953</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>368.5,-63.5,374.5,-63.5</points>
<intersection>368.5 0</intersection>
<intersection>374.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353.5,-114,353.5,-89</points>
<intersection>-114 1</intersection>
<intersection>-89 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326,-114,358,-114</points>
<connection>
<GID>952</GID>
<name>OUT_0</name></connection>
<connection>
<GID>954</GID>
<name>IN_1</name></connection>
<intersection>353.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>353.5,-89,359,-89</points>
<intersection>353.5 0</intersection>
<intersection>359 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>359,-97.5,359,-89</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<intersection>-89 4</intersection></vsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>340,-112,340,-96</points>
<intersection>-112 3</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325,-96,341.5,-96</points>
<connection>
<GID>950</GID>
<name>OUT_0</name></connection>
<intersection>340 0</intersection>
<intersection>341.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>340,-112,358,-112</points>
<connection>
<GID>954</GID>
<name>IN_0</name></connection>
<intersection>340 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>341.5,-96.5,341.5,-96</points>
<connection>
<GID>956</GID>
<name>IN_0</name></connection>
<intersection>-96 1</intersection></vsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-97.5,357,-96.5</points>
<connection>
<GID>958</GID>
<name>IN_1</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345.5,-96.5,357,-96.5</points>
<connection>
<GID>956</GID>
<name>OUT_0</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358,-104,363.5,-104</points>
<intersection>358 5</intersection>
<intersection>363.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>363.5,-104,363.5,-99.5</points>
<intersection>-104 1</intersection>
<intersection>-99.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>358,-104,358,-103.5</points>
<connection>
<GID>958</GID>
<name>OUT</name></connection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>363.5,-99.5,367,-99.5</points>
<connection>
<GID>1164</GID>
<name>IN_0</name></connection>
<intersection>363.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377.5,-99.5,377.5,-83</points>
<intersection>-99.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373,-99.5,377.5,-99.5</points>
<connection>
<GID>1164</GID>
<name>OUT_0</name></connection>
<intersection>377.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>377.5,-83,447,-83</points>
<connection>
<GID>1144</GID>
<name>IN_0</name></connection>
<intersection>377.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>373,-102.5,446,-102.5</points>
<connection>
<GID>1164</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>1146</GID>
<name>IN_1</name></connection>
<intersection>397.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>397.5,-207,397.5,-102.5</points>
<intersection>-207 8</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>397.5,-207,443,-207</points>
<connection>
<GID>970</GID>
<name>IN_3</name></connection>
<intersection>397.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>364,82.5,1007,82.5</points>
<intersection>364 15</intersection>
<intersection>371.5 16</intersection>
<intersection>1007 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>1007,-306,1007,82.5</points>
<intersection>-306 3</intersection>
<intersection>82.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>850,-306,1007,-306</points>
<intersection>850 14</intersection>
<intersection>866 13</intersection>
<intersection>879.5 12</intersection>
<intersection>894.5 11</intersection>
<intersection>905 10</intersection>
<intersection>918 9</intersection>
<intersection>1007 2</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>918,-306,918,-294.5</points>
<connection>
<GID>982</GID>
<name>clock</name></connection>
<intersection>-306 3</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>905,-306,905,-294.5</points>
<connection>
<GID>976</GID>
<name>clock</name></connection>
<intersection>-306 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>894.5,-306,894.5,-294.5</points>
<connection>
<GID>971</GID>
<name>clock</name></connection>
<intersection>-306 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>879.5,-306,879.5,-294.5</points>
<connection>
<GID>964</GID>
<name>clock</name></connection>
<intersection>-306 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>866,-306,866,-294.5</points>
<connection>
<GID>955</GID>
<name>clock</name></connection>
<intersection>-306 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>850,-306,850,-294</points>
<connection>
<GID>1145</GID>
<name>clock</name></connection>
<intersection>-306 3</intersection>
<intersection>-294 17</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>364,82.5,364,93</points>
<connection>
<GID>1034</GID>
<name>CLK</name></connection>
<intersection>82.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>371.5,82.5,371.5,93</points>
<connection>
<GID>1003</GID>
<name>IN_1</name></connection>
<intersection>82.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>767.5,-294,850,-294</points>
<intersection>767.5 18</intersection>
<intersection>850 14</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>767.5,-409,767.5,-294</points>
<intersection>-409 83</intersection>
<intersection>-294 17</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>849.5,-421,919,-421</points>
<intersection>849.5 52</intersection>
<intersection>867 51</intersection>
<intersection>880.5 50</intersection>
<intersection>895.5 49</intersection>
<intersection>906 48</intersection>
<intersection>919 47</intersection></hsegment>
<vsegment>
<ID>47</ID>
<points>919,-421,919,-409.5</points>
<connection>
<GID>1052</GID>
<name>clock</name></connection>
<intersection>-421 41</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>906,-421,906,-409.5</points>
<connection>
<GID>1050</GID>
<name>clock</name></connection>
<intersection>-421 41</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>895.5,-421,895.5,-409.5</points>
<connection>
<GID>1044</GID>
<name>clock</name></connection>
<intersection>-421 41</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>880.5,-421,880.5,-409.5</points>
<connection>
<GID>1039</GID>
<name>clock</name></connection>
<intersection>-421 41</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>867,-421,867,-409.5</points>
<connection>
<GID>1025</GID>
<name>clock</name></connection>
<intersection>-421 41</intersection></vsegment>
<vsegment>
<ID>52</ID>
<points>849.5,-421,849.5,-409</points>
<intersection>-421 41</intersection>
<intersection>-409 83</intersection></vsegment>
<hsegment>
<ID>83</ID>
<points>767.5,-409,851,-409</points>
<connection>
<GID>1124</GID>
<name>clock</name></connection>
<intersection>767.5 18</intersection>
<intersection>849.5 52</intersection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619.5,29.5,619.5,30.5</points>
<intersection>29.5 2</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>615,30.5,619.5,30.5</points>
<connection>
<GID>1001</GID>
<name>IN_1</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>619.5,29.5,624.5,29.5</points>
<connection>
<GID>990</GID>
<name>Q</name></connection>
<intersection>619.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,42,388.5,46.5</points>
<intersection>42 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>385,42,388.5,42</points>
<connection>
<GID>1008</GID>
<name>IN_1</name></connection>
<intersection>388.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>388.5,46.5,392,46.5</points>
<connection>
<GID>1007</GID>
<name>OUT</name></connection>
<intersection>388.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>541,58.5,636,58.5</points>
<connection>
<GID>984</GID>
<name>OUT_0</name></connection>
<intersection>636 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>636,29.5,636,58.5</points>
<intersection>29.5 10</intersection>
<intersection>58.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>630.5,29.5,636,29.5</points>
<connection>
<GID>990</GID>
<name>J</name></connection>
<intersection>636 3</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>379,29.5,609,29.5</points>
<connection>
<GID>1033</GID>
<name>clear</name></connection>
<connection>
<GID>1027</GID>
<name>clear</name></connection>
<connection>
<GID>1024</GID>
<name>clear</name></connection>
<connection>
<GID>1022</GID>
<name>clear</name></connection>
<connection>
<GID>1035</GID>
<name>clear</name></connection>
<connection>
<GID>1001</GID>
<name>OUT</name></connection>
<intersection>379 6</intersection>
<intersection>515.5 4</intersection>
<intersection>561 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>561,29,561,29.5</points>
<connection>
<GID>1030</GID>
<name>clear</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>515.5,-6.5,515.5,29.5</points>
<intersection>-6.5 5</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>515.5,-6.5,606.5,-6.5</points>
<intersection>515.5 4</intersection>
<intersection>524.5 13</intersection>
<intersection>541 12</intersection>
<intersection>555.5 11</intersection>
<intersection>572.5 10</intersection>
<intersection>588.5 9</intersection>
<intersection>606.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>379,29.5,379,49.5</points>
<intersection>29.5 1</intersection>
<intersection>49.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>378.5,49.5,379,49.5</points>
<connection>
<GID>1011</GID>
<name>IN_0</name></connection>
<intersection>379 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>606.5,-6.5,606.5,-5.5</points>
<connection>
<GID>1059</GID>
<name>clear</name></connection>
<intersection>-6.5 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>588.5,-6.5,588.5,-5.5</points>
<connection>
<GID>1057</GID>
<name>clear</name></connection>
<intersection>-6.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>572.5,-6.5,572.5,-5.5</points>
<connection>
<GID>1056</GID>
<name>clear</name></connection>
<intersection>-6.5 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>555.5,-6.5,555.5,-5.5</points>
<connection>
<GID>1053</GID>
<name>clear</name></connection>
<intersection>-6.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>541,-6.5,541,-5.5</points>
<connection>
<GID>1051</GID>
<name>clear</name></connection>
<intersection>-6.5 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>524.5,-6.5,524.5,-5.5</points>
<connection>
<GID>1048</GID>
<name>clear</name></connection>
<intersection>-6.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>385,40,425,40</points>
<connection>
<GID>1008</GID>
<name>IN_0</name></connection>
<intersection>425 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>425,38,425,40</points>
<connection>
<GID>1005</GID>
<name>OUT</name></connection>
<intersection>40 1</intersection></vsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,50.5,366.5,54.5</points>
<intersection>50.5 2</intersection>
<intersection>54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,54.5,366.5,54.5</points>
<connection>
<GID>1014</GID>
<name>IN_1</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>366.5,50.5,372.5,50.5</points>
<connection>
<GID>1011</GID>
<name>OUT</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>612.5,33.5,612.5,116.5</points>
<intersection>33.5 2</intersection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516,116.5,612.5,116.5</points>
<connection>
<GID>997</GID>
<name>IN_0</name></connection>
<intersection>612.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>612.5,33.5,624.5,33.5</points>
<connection>
<GID>990</GID>
<name>nQ</name></connection>
<intersection>612.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>387,102.5,432.5,102.5</points>
<connection>
<GID>1012</GID>
<name>clear</name></connection>
<connection>
<GID>1010</GID>
<name>clear</name></connection>
<connection>
<GID>1009</GID>
<name>clear</name></connection>
<intersection>387 13</intersection>
<intersection>432.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>432.5,101.5,432.5,102.5</points>
<connection>
<GID>1015</GID>
<name>clear</name></connection>
<intersection>101.5 5</intersection>
<intersection>102.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432.5,101.5,514,101.5</points>
<connection>
<GID>1018</GID>
<name>clear</name></connection>
<connection>
<GID>1017</GID>
<name>clear</name></connection>
<intersection>432.5 4</intersection>
<intersection>495 12</intersection>
<intersection>514 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>514,94.5,514,101.5</points>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection>
<intersection>101.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>495,101.5,495,108.5</points>
<connection>
<GID>1019</GID>
<name>OUT</name></connection>
<intersection>101.5 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>387,67.5,387,102.5</points>
<intersection>67.5 14</intersection>
<intersection>102.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>387,67.5,478,67.5</points>
<connection>
<GID>1071</GID>
<name>clear</name></connection>
<connection>
<GID>1070</GID>
<name>clear</name></connection>
<connection>
<GID>1069</GID>
<name>clear</name></connection>
<connection>
<GID>1068</GID>
<name>clear</name></connection>
<connection>
<GID>1067</GID>
<name>clear</name></connection>
<connection>
<GID>1065</GID>
<name>clear</name></connection>
<intersection>387 13</intersection></hsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>483,121,516,121</points>
<intersection>483 3</intersection>
<intersection>516 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>483,117,483,121</points>
<intersection>117 5</intersection>
<intersection>121 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>516,118.5,516,121</points>
<connection>
<GID>997</GID>
<name>IN_1</name></connection>
<intersection>121 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>482,117,483,117</points>
<connection>
<GID>1054</GID>
<name>OUT</name></connection>
<intersection>483 3</intersection></hsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>614,44,614,46.5</points>
<intersection>44 2</intersection>
<intersection>46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>614,46.5,618,46.5</points>
<connection>
<GID>1002</GID>
<name>IN_0</name></connection>
<intersection>614 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>610.5,44,614,44</points>
<connection>
<GID>1047</GID>
<name>OUT</name></connection>
<intersection>614 0</intersection></hsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>631,33.5,631,46.5</points>
<intersection>33.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>630.5,33.5,631,33.5</points>
<connection>
<GID>990</GID>
<name>K</name></connection>
<intersection>631 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>624,46.5,631,46.5</points>
<connection>
<GID>1002</GID>
<name>OUT_0</name></connection>
<intersection>631 0</intersection></hsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>367.5,41,379,41</points>
<connection>
<GID>1023</GID>
<name>IN_0</name></connection>
<connection>
<GID>1008</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,42,361.5,52.5</points>
<connection>
<GID>1023</GID>
<name>OUT</name></connection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,52.5,361.5,52.5</points>
<connection>
<GID>1014</GID>
<name>IN_0</name></connection>
<intersection>361.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>346,53.5,354,53.5</points>
<connection>
<GID>1029</GID>
<name>N_in1</name></connection>
<connection>
<GID>1014</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,109.5,505.5,117.5</points>
<intersection>109.5 1</intersection>
<intersection>117.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,109.5,505.5,109.5</points>
<connection>
<GID>1019</GID>
<name>IN_1</name></connection>
<intersection>505.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>505.5,117.5,510,117.5</points>
<connection>
<GID>997</GID>
<name>OUT</name></connection>
<intersection>505.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,25,505.5,107.5</points>
<intersection>25 3</intersection>
<intersection>107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,107.5,505.5,107.5</points>
<connection>
<GID>1019</GID>
<name>IN_0</name></connection>
<intersection>505.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>366,25,615,25</points>
<connection>
<GID>1006</GID>
<name>OUT_0</name></connection>
<intersection>505.5 0</intersection>
<intersection>615 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>615,25,615,28.5</points>
<connection>
<GID>1001</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></vsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,104.5,412,117</points>
<intersection>104.5 4</intersection>
<intersection>108.5 2</intersection>
<intersection>117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>410.5,117,421.5,117</points>
<connection>
<GID>1037</GID>
<name>OUT</name></connection>
<connection>
<GID>1042</GID>
<name>IN_0</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412,108.5,413.5,108.5</points>
<connection>
<GID>1012</GID>
<name>J</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>412,104.5,413.5,104.5</points>
<connection>
<GID>1012</GID>
<name>K</name></connection>
<intersection>412 0</intersection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,104,428.5,116</points>
<intersection>104 4</intersection>
<intersection>108 2</intersection>
<intersection>116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,116,436.5,116</points>
<connection>
<GID>1042</GID>
<name>OUT</name></connection>
<connection>
<GID>1046</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>428.5,108,429.5,108</points>
<connection>
<GID>1015</GID>
<name>J</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>428.5,104,429.5,104</points>
<connection>
<GID>1015</GID>
<name>K</name></connection>
<intersection>428.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,103.5,444,115</points>
<intersection>103.5 4</intersection>
<intersection>107.5 2</intersection>
<intersection>115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,115,454,115</points>
<connection>
<GID>1046</GID>
<name>OUT</name></connection>
<connection>
<GID>1049</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,107.5,445.5,107.5</points>
<connection>
<GID>1017</GID>
<name>J</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>444,103.5,445.5,103.5</points>
<connection>
<GID>1017</GID>
<name>K</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461,103.5,461,114</points>
<intersection>103.5 4</intersection>
<intersection>107.5 2</intersection>
<intersection>114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>460,114,461,114</points>
<connection>
<GID>1049</GID>
<name>OUT</name></connection>
<intersection>461 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>461,107.5,462.5,107.5</points>
<connection>
<GID>1018</GID>
<name>J</name></connection>
<intersection>461 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>461,103.5,462.5,103.5</points>
<connection>
<GID>1018</GID>
<name>K</name></connection>
<intersection>461 0</intersection></hsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>390,108.5,397.5,108.5</points>
<connection>
<GID>1009</GID>
<name>Q</name></connection>
<connection>
<GID>1010</GID>
<name>J</name></connection>
<intersection>391 3</intersection>
<intersection>393.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>391,73.5,391,108.5</points>
<intersection>73.5 10</intersection>
<intersection>89 4</intersection>
<intersection>104.5 9</intersection>
<intersection>108.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>391,89,478,89</points>
<connection>
<GID>1026</GID>
<name>IN_0</name></connection>
<intersection>391 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>393.5,108.5,393.5,118</points>
<intersection>108.5 1</intersection>
<intersection>118 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>393.5,118,404.5,118</points>
<connection>
<GID>1037</GID>
<name>IN_0</name></connection>
<intersection>393.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>391,104.5,397.5,104.5</points>
<connection>
<GID>1010</GID>
<name>K</name></connection>
<intersection>391 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>391,73.5,393,73.5</points>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection>
<intersection>391 3</intersection></hsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>378,99,632.5,99</points>
<intersection>378 3</intersection>
<intersection>393.5 4</intersection>
<intersection>409.5 32</intersection>
<intersection>410.5 5</intersection>
<intersection>424 31</intersection>
<intersection>426.5 16</intersection>
<intersection>441 30</intersection>
<intersection>443 15</intersection>
<intersection>457 29</intersection>
<intersection>458 18</intersection>
<intersection>475 28</intersection>
<intersection>632.5 35</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>378,70.5,378,106.5</points>
<intersection>70.5 33</intersection>
<intersection>94 39</intersection>
<intersection>99 1</intersection>
<intersection>106.5 13</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>393.5,99,393.5,106.5</points>
<intersection>99 1</intersection>
<intersection>106.5 14</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>410.5,99,410.5,106.5</points>
<intersection>99 1</intersection>
<intersection>106.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>410.5,106.5,413.5,106.5</points>
<connection>
<GID>1012</GID>
<name>clock</name></connection>
<intersection>410.5 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>378,106.5,384,106.5</points>
<connection>
<GID>1009</GID>
<name>clock</name></connection>
<intersection>378 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>393.5,106.5,397.5,106.5</points>
<connection>
<GID>1010</GID>
<name>clock</name></connection>
<intersection>393.5 4</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>443,99,443,105.5</points>
<intersection>99 1</intersection>
<intersection>105.5 21</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>426.5,99,426.5,106</points>
<intersection>99 1</intersection>
<intersection>106 19</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>458,99,458,105.5</points>
<intersection>99 1</intersection>
<intersection>105.5 20</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>426.5,106,429.5,106</points>
<connection>
<GID>1015</GID>
<name>clock</name></connection>
<intersection>426.5 16</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>458,105.5,462.5,105.5</points>
<connection>
<GID>1018</GID>
<name>clock</name></connection>
<intersection>458 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>443,105.5,445.5,105.5</points>
<connection>
<GID>1017</GID>
<name>clock</name></connection>
<intersection>443 15</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>475,70.5,475,99</points>
<connection>
<GID>1071</GID>
<name>clock</name></connection>
<intersection>99 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>457,70.5,457,99</points>
<connection>
<GID>1070</GID>
<name>clock</name></connection>
<intersection>99 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>441,70.5,441,99</points>
<connection>
<GID>1069</GID>
<name>clock</name></connection>
<intersection>99 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>424,70.5,424,99</points>
<connection>
<GID>1068</GID>
<name>clock</name></connection>
<intersection>99 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>409.5,70.5,409.5,99</points>
<connection>
<GID>1067</GID>
<name>clock</name></connection>
<intersection>99 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>378,70.5,393,70.5</points>
<connection>
<GID>1065</GID>
<name>clock</name></connection>
<intersection>378 3</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>632.5,31.5,632.5,99</points>
<intersection>31.5 36</intersection>
<intersection>99 1</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>630.5,31.5,632.5,31.5</points>
<connection>
<GID>990</GID>
<name>clock</name></connection>
<intersection>632.5 35</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>377.5,94,378,94</points>
<connection>
<GID>1003</GID>
<name>OUT</name></connection>
<intersection>378 3</intersection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404.5,73.5,404.5,116</points>
<connection>
<GID>1037</GID>
<name>IN_1</name></connection>
<intersection>73.5 8</intersection>
<intersection>90 1</intersection>
<intersection>108.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>404.5,90,478,90</points>
<connection>
<GID>1026</GID>
<name>IN_1</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>403.5,108.5,404.5,108.5</points>
<connection>
<GID>1010</GID>
<name>Q</name></connection>
<intersection>404.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>404.5,73.5,409.5,73.5</points>
<connection>
<GID>1067</GID>
<name>IN_0</name></connection>
<intersection>404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>436.5,92,478,92</points>
<connection>
<GID>1026</GID>
<name>IN_3</name></connection>
<intersection>436.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>436.5,73.5,436.5,118</points>
<connection>
<GID>1046</GID>
<name>IN_1</name></connection>
<intersection>73.5 9</intersection>
<intersection>92 1</intersection>
<intersection>108 4</intersection>
<intersection>118 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>435.5,108,436.5,108</points>
<connection>
<GID>1015</GID>
<name>Q</name></connection>
<intersection>436.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>436.5,118,476,118</points>
<connection>
<GID>1054</GID>
<name>IN_1</name></connection>
<intersection>436.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>436.5,73.5,441,73.5</points>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection>
<intersection>436.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420.5,73.5,420.5,120</points>
<intersection>73.5 9</intersection>
<intersection>91 4</intersection>
<intersection>108.5 3</intersection>
<intersection>115 2</intersection>
<intersection>120 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>420.5,115,421.5,115</points>
<connection>
<GID>1042</GID>
<name>IN_1</name></connection>
<intersection>420.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>419.5,108.5,420.5,108.5</points>
<connection>
<GID>1012</GID>
<name>Q</name></connection>
<intersection>420.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>420.5,91,478,91</points>
<connection>
<GID>1026</GID>
<name>IN_2</name></connection>
<intersection>420.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>420.5,120,476,120</points>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection>
<intersection>420.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>420.5,73.5,424,73.5</points>
<connection>
<GID>1068</GID>
<name>IN_0</name></connection>
<intersection>420.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,73.5,452.5,116</points>
<intersection>73.5 8</intersection>
<intersection>93 3</intersection>
<intersection>107.5 1</intersection>
<intersection>116 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>451.5,107.5,452.5,107.5</points>
<connection>
<GID>1017</GID>
<name>Q</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>452.5,116,476,116</points>
<connection>
<GID>1054</GID>
<name>IN_2</name></connection>
<intersection>452.5 0</intersection>
<intersection>454 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>452.5,93,478,93</points>
<connection>
<GID>1026</GID>
<name>IN_4</name></connection>
<intersection>452.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>454,113,454,116</points>
<connection>
<GID>1049</GID>
<name>IN_1</name></connection>
<intersection>116 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>452.5,73.5,457,73.5</points>
<connection>
<GID>1070</GID>
<name>IN_0</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470.5,73.5,470.5,114</points>
<intersection>73.5 5</intersection>
<intersection>94 2</intersection>
<intersection>107.5 1</intersection>
<intersection>114 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>468.5,107.5,470.5,107.5</points>
<connection>
<GID>1018</GID>
<name>Q</name></connection>
<intersection>470.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>470.5,94,478,94</points>
<connection>
<GID>1026</GID>
<name>IN_5</name></connection>
<intersection>470.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>470.5,114,476,114</points>
<connection>
<GID>1054</GID>
<name>IN_3</name></connection>
<intersection>470.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>470.5,73.5,475,73.5</points>
<connection>
<GID>1071</GID>
<name>IN_0</name></connection>
<intersection>470.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>400.5,59,493,59</points>
<connection>
<GID>1072</GID>
<name>IN_0</name></connection>
<intersection>400.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>400.5,49.5,400.5,73.5</points>
<intersection>49.5 8</intersection>
<intersection>59 1</intersection>
<intersection>73.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>399,73.5,400.5,73.5</points>
<connection>
<GID>1065</GID>
<name>OUT_0</name></connection>
<intersection>400.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>399,49.5,400.5,49.5</points>
<connection>
<GID>1007</GID>
<name>IN_3</name></connection>
<intersection>400.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>417,60,493,60</points>
<connection>
<GID>1072</GID>
<name>IN_1</name></connection>
<intersection>417 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>417,47.5,417,73.5</points>
<intersection>47.5 8</intersection>
<intersection>60 1</intersection>
<intersection>73.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>415.5,73.5,417,73.5</points>
<connection>
<GID>1067</GID>
<name>OUT_0</name></connection>
<intersection>417 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>399,47.5,417,47.5</points>
<connection>
<GID>1007</GID>
<name>IN_2</name></connection>
<intersection>417 3</intersection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431,61,493,61</points>
<connection>
<GID>1072</GID>
<name>IN_2</name></connection>
<intersection>431 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>431,45.5,431,73.5</points>
<intersection>45.5 8</intersection>
<intersection>61 1</intersection>
<intersection>73.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>430,73.5,431,73.5</points>
<connection>
<GID>1068</GID>
<name>OUT_0</name></connection>
<intersection>431 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>399,45.5,431,45.5</points>
<connection>
<GID>1007</GID>
<name>IN_1</name></connection>
<intersection>431 3</intersection></hsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449.5,62,493,62</points>
<connection>
<GID>1072</GID>
<name>IN_3</name></connection>
<intersection>449.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449.5,43.5,449.5,73.5</points>
<intersection>43.5 8</intersection>
<intersection>62 1</intersection>
<intersection>73.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>447,73.5,449.5,73.5</points>
<connection>
<GID>1069</GID>
<name>OUT_0</name></connection>
<intersection>449.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>399,43.5,449.5,43.5</points>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection>
<intersection>449.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>431,63,493,63</points>
<connection>
<GID>1072</GID>
<name>IN_4</name></connection>
<intersection>431 7</intersection>
<intersection>464 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>464,63,464,73.5</points>
<intersection>63 1</intersection>
<intersection>73.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>463,73.5,464,73.5</points>
<connection>
<GID>1070</GID>
<name>OUT_0</name></connection>
<intersection>464 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>431,39,431,63</points>
<connection>
<GID>1005</GID>
<name>IN_1</name></connection>
<intersection>63 1</intersection></vsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>484,64,493,64</points>
<connection>
<GID>1072</GID>
<name>IN_5</name></connection>
<intersection>484 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>484,37,484,73.5</points>
<intersection>37 8</intersection>
<intersection>64 1</intersection>
<intersection>73.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>481,73.5,484,73.5</points>
<connection>
<GID>1071</GID>
<name>OUT_0</name></connection>
<intersection>484 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>431,37,484,37</points>
<connection>
<GID>1005</GID>
<name>IN_0</name></connection>
<intersection>484 5</intersection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,31.5,540.5,44</points>
<intersection>31.5 4</intersection>
<intersection>35.5 2</intersection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>539,44,550,44</points>
<connection>
<GID>1040</GID>
<name>OUT</name></connection>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,35.5,542,35.5</points>
<connection>
<GID>1027</GID>
<name>J</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>540.5,31.5,542,31.5</points>
<connection>
<GID>1027</GID>
<name>K</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>557,31,557,43</points>
<intersection>31 4</intersection>
<intersection>35 2</intersection>
<intersection>43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>556,43,565,43</points>
<connection>
<GID>1041</GID>
<name>OUT</name></connection>
<connection>
<GID>1043</GID>
<name>IN_0</name></connection>
<intersection>557 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>557,35,558,35</points>
<connection>
<GID>1030</GID>
<name>J</name></connection>
<intersection>557 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>557,31,558,31</points>
<connection>
<GID>1030</GID>
<name>K</name></connection>
<intersection>557 0</intersection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572.5,31.5,572.5,42</points>
<intersection>31.5 4</intersection>
<intersection>35.5 2</intersection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571,42,582.5,42</points>
<connection>
<GID>1043</GID>
<name>OUT</name></connection>
<connection>
<GID>1045</GID>
<name>IN_0</name></connection>
<intersection>572.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>572.5,35.5,574,35.5</points>
<connection>
<GID>1033</GID>
<name>J</name></connection>
<intersection>572.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>572.5,31.5,574,31.5</points>
<connection>
<GID>1033</GID>
<name>K</name></connection>
<intersection>572.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,31.5,589.5,41</points>
<intersection>31.5 4</intersection>
<intersection>35.5 2</intersection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>588.5,41,589.5,41</points>
<connection>
<GID>1045</GID>
<name>OUT</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,35.5,591,35.5</points>
<connection>
<GID>1035</GID>
<name>J</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>589.5,31.5,591,31.5</points>
<connection>
<GID>1035</GID>
<name>K</name></connection>
<intersection>589.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>518.5,35.5,526,35.5</points>
<connection>
<GID>1022</GID>
<name>Q</name></connection>
<connection>
<GID>1024</GID>
<name>J</name></connection>
<intersection>519.5 3</intersection>
<intersection>522 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>519.5,0.5,519.5,35.5</points>
<intersection>0.5 10</intersection>
<intersection>16 4</intersection>
<intersection>31.5 9</intersection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>519.5,16,601,16</points>
<connection>
<GID>1036</GID>
<name>IN_0</name></connection>
<intersection>519.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>522,35.5,522,45</points>
<intersection>35.5 1</intersection>
<intersection>45 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>522,45,533,45</points>
<connection>
<GID>1040</GID>
<name>IN_0</name></connection>
<intersection>522 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>519.5,31.5,526,31.5</points>
<connection>
<GID>1024</GID>
<name>K</name></connection>
<intersection>519.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>519.5,0.5,521.5,0.5</points>
<connection>
<GID>1048</GID>
<name>IN_0</name></connection>
<intersection>519.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,0.5,533,43</points>
<connection>
<GID>1040</GID>
<name>IN_1</name></connection>
<intersection>0.5 8</intersection>
<intersection>17 1</intersection>
<intersection>35.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>533,17,601,17</points>
<connection>
<GID>1036</GID>
<name>IN_1</name></connection>
<intersection>533 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>532,35.5,533,35.5</points>
<connection>
<GID>1024</GID>
<name>Q</name></connection>
<intersection>533 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>533,0.5,538,0.5</points>
<connection>
<GID>1051</GID>
<name>IN_0</name></connection>
<intersection>533 0</intersection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>565,19,601,19</points>
<connection>
<GID>1036</GID>
<name>IN_3</name></connection>
<intersection>565 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>565,0.5,565,45</points>
<connection>
<GID>1043</GID>
<name>IN_1</name></connection>
<intersection>0.5 9</intersection>
<intersection>19 1</intersection>
<intersection>35 4</intersection>
<intersection>45 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>564,35,565,35</points>
<connection>
<GID>1030</GID>
<name>Q</name></connection>
<intersection>565 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>565,45,604.5,45</points>
<connection>
<GID>1047</GID>
<name>IN_1</name></connection>
<intersection>565 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>565,0.5,569.5,0.5</points>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection>
<intersection>565 3</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>549,0.5,549,47</points>
<intersection>0.5 9</intersection>
<intersection>18 4</intersection>
<intersection>35.5 3</intersection>
<intersection>42 2</intersection>
<intersection>47 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>549,42,550,42</points>
<connection>
<GID>1041</GID>
<name>IN_1</name></connection>
<intersection>549 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>548,35.5,549,35.5</points>
<connection>
<GID>1027</GID>
<name>Q</name></connection>
<intersection>549 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>549,18,601,18</points>
<connection>
<GID>1036</GID>
<name>IN_2</name></connection>
<intersection>549 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>549,47,604.5,47</points>
<connection>
<GID>1047</GID>
<name>IN_0</name></connection>
<intersection>549 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>549,0.5,552.5,0.5</points>
<connection>
<GID>1053</GID>
<name>IN_0</name></connection>
<intersection>549 0</intersection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,0.5,581,43</points>
<intersection>0.5 8</intersection>
<intersection>20 3</intersection>
<intersection>35.5 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>580,35.5,581,35.5</points>
<connection>
<GID>1033</GID>
<name>Q</name></connection>
<intersection>581 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>581,43,604.5,43</points>
<connection>
<GID>1047</GID>
<name>IN_2</name></connection>
<intersection>581 0</intersection>
<intersection>582.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>581,20,601,20</points>
<connection>
<GID>1036</GID>
<name>IN_4</name></connection>
<intersection>581 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>582.5,40,582.5,43</points>
<connection>
<GID>1045</GID>
<name>IN_1</name></connection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>581,0.5,585.5,0.5</points>
<connection>
<GID>1057</GID>
<name>IN_0</name></connection>
<intersection>581 0</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>599,0.5,599,41</points>
<intersection>0.5 5</intersection>
<intersection>21 2</intersection>
<intersection>35.5 1</intersection>
<intersection>41 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597,35.5,599,35.5</points>
<connection>
<GID>1035</GID>
<name>Q</name></connection>
<intersection>599 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>599,21,601,21</points>
<connection>
<GID>1036</GID>
<name>IN_5</name></connection>
<intersection>599 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>599,41,604.5,41</points>
<connection>
<GID>1047</GID>
<name>IN_3</name></connection>
<intersection>599 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>599,0.5,603.5,0.5</points>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection>
<intersection>599 0</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>529,-51.5,842.5,-51.5</points>
<intersection>529 3</intersection>
<intersection>842.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>529,-51.5,529,0.5</points>
<intersection>-51.5 1</intersection>
<intersection>-14 7</intersection>
<intersection>0.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>527.5,0.5,529,0.5</points>
<connection>
<GID>1048</GID>
<name>OUT_0</name></connection>
<intersection>529 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>842.5,-320,842.5,-51.5</points>
<intersection>-320 10</intersection>
<intersection>-278.5 11</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>529,-14,621.5,-14</points>
<connection>
<GID>1061</GID>
<name>IN_0</name></connection>
<intersection>529 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>842.5,-320,851,-320</points>
<intersection>842.5 5</intersection>
<intersection>851 12</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>842.5,-278.5,850,-278.5</points>
<intersection>842.5 5</intersection>
<intersection>850 13</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>851,-396.5,851,-320</points>
<connection>
<GID>1118</GID>
<name>IN_0</name></connection>
<intersection>-320 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>850,-281.5,850,-278.5</points>
<connection>
<GID>1076</GID>
<name>IN_0</name></connection>
<intersection>-278.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>545.5,-47,864.5,-47</points>
<intersection>545.5 3</intersection>
<intersection>864.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>545.5,-47,545.5,0.5</points>
<intersection>-47 1</intersection>
<intersection>-13 7</intersection>
<intersection>0.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>544,0.5,545.5,0.5</points>
<connection>
<GID>1051</GID>
<name>OUT_0</name></connection>
<intersection>545.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>864.5,-396.5,864.5,-47</points>
<connection>
<GID>1119</GID>
<name>IN_0</name></connection>
<intersection>-281.5 9</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>545.5,-13,621.5,-13</points>
<connection>
<GID>1061</GID>
<name>IN_1</name></connection>
<intersection>545.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>863.5,-281.5,864.5,-281.5</points>
<connection>
<GID>1077</GID>
<name>IN_0</name></connection>
<intersection>864.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>559.5,-42.5,877.5,-42.5</points>
<intersection>559.5 3</intersection>
<intersection>877.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>559.5,-42.5,559.5,0.5</points>
<intersection>-42.5 1</intersection>
<intersection>-12 7</intersection>
<intersection>0.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>558.5,0.5,559.5,0.5</points>
<connection>
<GID>1053</GID>
<name>OUT_0</name></connection>
<intersection>559.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>877.5,-396.5,877.5,-42.5</points>
<connection>
<GID>1120</GID>
<name>IN_0</name></connection>
<intersection>-281.5 9</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>559.5,-12,621.5,-12</points>
<connection>
<GID>1061</GID>
<name>IN_2</name></connection>
<intersection>559.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>876.5,-281.5,877.5,-281.5</points>
<connection>
<GID>1079</GID>
<name>IN_0</name></connection>
<intersection>877.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578,-38,890.5,-38</points>
<intersection>578 3</intersection>
<intersection>890.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>578,-38,578,0.5</points>
<intersection>-38 1</intersection>
<intersection>-11 7</intersection>
<intersection>0.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>575.5,0.5,578,0.5</points>
<connection>
<GID>1056</GID>
<name>OUT_0</name></connection>
<intersection>578 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>890.5,-396.5,890.5,-38</points>
<connection>
<GID>1121</GID>
<name>IN_0</name></connection>
<intersection>-281.5 9</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>578,-11,621.5,-11</points>
<connection>
<GID>1061</GID>
<name>IN_3</name></connection>
<intersection>578 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>889.5,-281.5,890.5,-281.5</points>
<connection>
<GID>1081</GID>
<name>IN_0</name></connection>
<intersection>890.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593,-35,903,-35</points>
<intersection>593 3</intersection>
<intersection>903 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>593,-35,593,0.5</points>
<intersection>-35 1</intersection>
<intersection>-10 7</intersection>
<intersection>0.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>591.5,0.5,593,0.5</points>
<connection>
<GID>1057</GID>
<name>OUT_0</name></connection>
<intersection>593 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>903,-397,903,-35</points>
<connection>
<GID>1122</GID>
<name>IN_0</name></connection>
<intersection>-282 9</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>593,-10,621.5,-10</points>
<connection>
<GID>1061</GID>
<name>IN_4</name></connection>
<intersection>593 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>902,-282,903,-282</points>
<connection>
<GID>1082</GID>
<name>IN_0</name></connection>
<intersection>903 5</intersection></hsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>615.5,-30,615.5,0.5</points>
<intersection>-30 5</intersection>
<intersection>-9 8</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>609.5,0.5,615.5,0.5</points>
<connection>
<GID>1059</GID>
<name>OUT_0</name></connection>
<intersection>615.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>615.5,-30,915.5,-30</points>
<intersection>615.5 0</intersection>
<intersection>915.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>915.5,-397,915.5,-30</points>
<connection>
<GID>1123</GID>
<name>IN_0</name></connection>
<intersection>-282 10</intersection>
<intersection>-30 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>615.5,-9,621.5,-9</points>
<connection>
<GID>1061</GID>
<name>IN_5</name></connection>
<intersection>615.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>914.5,-282,915.5,-282</points>
<connection>
<GID>1084</GID>
<name>IN_0</name></connection>
<intersection>915.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>509,31.5,509,58.5</points>
<intersection>31.5 4</intersection>
<intersection>35.5 17</intersection>
<intersection>58.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>370,31.5,512.5,31.5</points>
<connection>
<GID>1022</GID>
<name>K</name></connection>
<intersection>370 11</intersection>
<intersection>509 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>509,58.5,535,58.5</points>
<connection>
<GID>984</GID>
<name>IN_0</name></connection>
<intersection>509 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>370,108.5,384,108.5</points>
<connection>
<GID>1009</GID>
<name>J</name></connection>
<intersection>370 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>370,31.5,370,108.5</points>
<intersection>31.5 4</intersection>
<intersection>43 22</intersection>
<intersection>56 23</intersection>
<intersection>95 21</intersection>
<intersection>102.5 28</intersection>
<intersection>104.5 14</intersection>
<intersection>108.5 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>370,104.5,384,104.5</points>
<connection>
<GID>1009</GID>
<name>K</name></connection>
<intersection>370 11</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>509,35.5,512.5,35.5</points>
<connection>
<GID>1022</GID>
<name>J</name></connection>
<intersection>509 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>370,95,371.5,95</points>
<connection>
<GID>1003</GID>
<name>IN_0</name></connection>
<intersection>370 11</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>367.5,43,370,43</points>
<connection>
<GID>1023</GID>
<name>IN_1</name></connection>
<intersection>370 11</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>370,56,378.5,56</points>
<intersection>370 11</intersection>
<intersection>378.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>378.5,51.5,378.5,56</points>
<connection>
<GID>1011</GID>
<name>IN_1</name></connection>
<intersection>56 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>363.5,102.5,370,102.5</points>
<connection>
<GID>1073</GID>
<name>OUT</name></connection>
<intersection>370 11</intersection></hsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-2.5,511.5,88.5</points>
<intersection>-2.5 8</intersection>
<intersection>33.5 1</intersection>
<intersection>88.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511.5,33.5,591,33.5</points>
<connection>
<GID>1022</GID>
<name>clock</name></connection>
<connection>
<GID>1024</GID>
<name>clock</name></connection>
<connection>
<GID>1027</GID>
<name>clock</name></connection>
<connection>
<GID>1033</GID>
<name>clock</name></connection>
<connection>
<GID>1035</GID>
<name>clock</name></connection>
<intersection>511.5 0</intersection>
<intersection>558 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>558,33,558,33.5</points>
<connection>
<GID>1030</GID>
<name>clock</name></connection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>511.5,-2.5,603.5,-2.5</points>
<connection>
<GID>1048</GID>
<name>clock</name></connection>
<connection>
<GID>1051</GID>
<name>clock</name></connection>
<connection>
<GID>1053</GID>
<name>clock</name></connection>
<connection>
<GID>1056</GID>
<name>clock</name></connection>
<connection>
<GID>1057</GID>
<name>clock</name></connection>
<connection>
<GID>1059</GID>
<name>clock</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>511.5,88.5,514,88.5</points>
<connection>
<GID>1063</GID>
<name>OUT_0</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>735.5,-391,735.5,-333</points>
<connection>
<GID>1088</GID>
<name>OUT_0</name></connection>
<intersection>-391 1</intersection>
<intersection>-382.5 7</intersection>
<intersection>-374 3</intersection>
<intersection>-366 8</intersection>
<intersection>-357.5 5</intersection>
<intersection>-349 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>735.5,-391,758.5,-391</points>
<connection>
<GID>1089</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>735.5,-374,757.5,-374</points>
<connection>
<GID>1091</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>735.5,-357.5,756.5,-357.5</points>
<connection>
<GID>1093</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>735.5,-382.5,758,-382.5</points>
<connection>
<GID>1090</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>735.5,-366,757,-366</points>
<connection>
<GID>1092</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>735.5,-349,756.5,-349</points>
<connection>
<GID>1094</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>894.5,-452.5,894.5,-447.5</points>
<connection>
<GID>1117</GID>
<name>OUT</name></connection>
<intersection>-452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>894.5,-452.5,911,-452.5</points>
<connection>
<GID>1097</GID>
<name>N_in0</name></connection>
<intersection>894.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>766,-245.5,825,-245.5</points>
<connection>
<GID>1125</GID>
<name>OUT</name></connection>
<connection>
<GID>1098</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>848,-281.5,848,-245.5</points>
<connection>
<GID>1076</GID>
<name>IN_1</name></connection>
<intersection>-245.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>831,-245.5,848,-245.5</points>
<connection>
<GID>1098</GID>
<name>Q</name></connection>
<intersection>848 0</intersection></hsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>765.5,-235.5,812,-235.5</points>
<connection>
<GID>1126</GID>
<name>OUT</name></connection>
<connection>
<GID>1099</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>861.5,-281.5,861.5,-235.5</points>
<connection>
<GID>1077</GID>
<name>IN_1</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>818,-235.5,861.5,-235.5</points>
<connection>
<GID>1099</GID>
<name>Q</name></connection>
<intersection>861.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>764,-224.5,799,-224.5</points>
<connection>
<GID>1127</GID>
<name>OUT</name></connection>
<connection>
<GID>1100</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>874.5,-281.5,874.5,-224.5</points>
<connection>
<GID>1079</GID>
<name>IN_1</name></connection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>805,-224.5,874.5,-224.5</points>
<connection>
<GID>1100</GID>
<name>Q</name></connection>
<intersection>874.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>763.5,-215.5,791.5,-215.5</points>
<connection>
<GID>1128</GID>
<name>OUT</name></connection>
<connection>
<GID>1101</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>887.5,-281.5,887.5,-215.5</points>
<connection>
<GID>1081</GID>
<name>IN_1</name></connection>
<intersection>-215.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>797.5,-215.5,887.5,-215.5</points>
<connection>
<GID>1101</GID>
<name>Q</name></connection>
<intersection>887.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>762.5,-208,783,-208</points>
<connection>
<GID>1129</GID>
<name>OUT</name></connection>
<connection>
<GID>1102</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>900,-282,900,-208</points>
<connection>
<GID>1082</GID>
<name>IN_1</name></connection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>789,-208,900,-208</points>
<connection>
<GID>1102</GID>
<name>Q</name></connection>
<intersection>900 0</intersection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>761.5,-200.5,774,-200.5</points>
<connection>
<GID>1130</GID>
<name>OUT</name></connection>
<connection>
<GID>1103</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>912.5,-282,912.5,-200.5</points>
<connection>
<GID>1084</GID>
<name>IN_1</name></connection>
<intersection>-200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>780,-200.5,912.5,-200.5</points>
<connection>
<GID>1103</GID>
<name>Q</name></connection>
<intersection>912.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>764.5,-392,816.5,-392</points>
<connection>
<GID>1089</GID>
<name>OUT</name></connection>
<connection>
<GID>1104</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>849,-396.5,849,-392</points>
<connection>
<GID>1118</GID>
<name>IN_1</name></connection>
<intersection>-392 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>822.5,-392,849,-392</points>
<connection>
<GID>1104</GID>
<name>Q</name></connection>
<intersection>849 0</intersection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>764,-383.5,808.5,-383.5</points>
<connection>
<GID>1090</GID>
<name>OUT</name></connection>
<connection>
<GID>1105</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>862.5,-396.5,862.5,-383.5</points>
<connection>
<GID>1119</GID>
<name>IN_1</name></connection>
<intersection>-383.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>814.5,-383.5,862.5,-383.5</points>
<connection>
<GID>1105</GID>
<name>Q</name></connection>
<intersection>862.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>763.5,-375,801.5,-375</points>
<connection>
<GID>1091</GID>
<name>OUT</name></connection>
<connection>
<GID>1106</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>875.5,-396.5,875.5,-375</points>
<connection>
<GID>1120</GID>
<name>IN_1</name></connection>
<intersection>-375 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>807.5,-375,875.5,-375</points>
<connection>
<GID>1106</GID>
<name>Q</name></connection>
<intersection>875.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>763,-367,792.5,-367</points>
<connection>
<GID>1092</GID>
<name>OUT</name></connection>
<connection>
<GID>1107</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>888.5,-396.5,888.5,-367</points>
<connection>
<GID>1121</GID>
<name>IN_1</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>798.5,-367,888.5,-367</points>
<connection>
<GID>1107</GID>
<name>Q</name></connection>
<intersection>888.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>762.5,-358.5,785.5,-358.5</points>
<connection>
<GID>1093</GID>
<name>OUT</name></connection>
<connection>
<GID>1108</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>901,-397,901,-358.5</points>
<connection>
<GID>1122</GID>
<name>IN_1</name></connection>
<intersection>-358.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>791.5,-358.5,901,-358.5</points>
<connection>
<GID>1108</GID>
<name>Q</name></connection>
<intersection>901 0</intersection></hsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>762.5,-350,777.5,-350</points>
<connection>
<GID>1094</GID>
<name>OUT</name></connection>
<connection>
<GID>1109</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>913.5,-397,913.5,-350</points>
<connection>
<GID>1123</GID>
<name>IN_1</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>783.5,-350,913.5,-350</points>
<connection>
<GID>1109</GID>
<name>Q</name></connection>
<intersection>913.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>780.5,-398,780.5,-356</points>
<connection>
<GID>1109</GID>
<name>clear</name></connection>
<intersection>-398 10</intersection>
<intersection>-389.5 5</intersection>
<intersection>-381 9</intersection>
<intersection>-373 3</intersection>
<intersection>-364.5 7</intersection>
<intersection>-356 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>780.5,-356,808.5,-356</points>
<connection>
<GID>1110</GID>
<name>OUT_0</name></connection>
<intersection>780.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>780.5,-373,795.5,-373</points>
<connection>
<GID>1107</GID>
<name>clear</name></connection>
<intersection>780.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>780.5,-389.5,811.5,-389.5</points>
<connection>
<GID>1105</GID>
<name>clear</name></connection>
<intersection>780.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>780.5,-364.5,788.5,-364.5</points>
<connection>
<GID>1108</GID>
<name>clear</name></connection>
<intersection>780.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>780.5,-381,804.5,-381</points>
<connection>
<GID>1106</GID>
<name>clear</name></connection>
<intersection>780.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>780.5,-398,819.5,-398</points>
<connection>
<GID>1104</GID>
<name>clear</name></connection>
<intersection>780.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>773,-394,773,-346</points>
<connection>
<GID>1112</GID>
<name>OUT_0</name></connection>
<intersection>-394 7</intersection>
<intersection>-385.5 5</intersection>
<intersection>-377 8</intersection>
<intersection>-369 3</intersection>
<intersection>-360.5 9</intersection>
<intersection>-352 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>773,-352,777.5,-352</points>
<connection>
<GID>1109</GID>
<name>clock</name></connection>
<intersection>773 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>773,-369,792.5,-369</points>
<connection>
<GID>1107</GID>
<name>clock</name></connection>
<intersection>773 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>773,-385.5,808.5,-385.5</points>
<connection>
<GID>1105</GID>
<name>clock</name></connection>
<intersection>773 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>773,-394,816.5,-394</points>
<connection>
<GID>1104</GID>
<name>clock</name></connection>
<intersection>773 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>773,-377,801.5,-377</points>
<connection>
<GID>1106</GID>
<name>clock</name></connection>
<intersection>773 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>773,-360.5,785.5,-360.5</points>
<connection>
<GID>1108</GID>
<name>clock</name></connection>
<intersection>773 0</intersection></hsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>769.5,-247.5,769.5,-196.5</points>
<connection>
<GID>1113</GID>
<name>OUT_0</name></connection>
<intersection>-247.5 7</intersection>
<intersection>-237.5 5</intersection>
<intersection>-226.5 8</intersection>
<intersection>-217.5 3</intersection>
<intersection>-210 9</intersection>
<intersection>-202.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>769.5,-202.5,774,-202.5</points>
<connection>
<GID>1103</GID>
<name>clock</name></connection>
<intersection>769.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>769.5,-217.5,791.5,-217.5</points>
<connection>
<GID>1101</GID>
<name>clock</name></connection>
<intersection>769.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>769.5,-237.5,812,-237.5</points>
<connection>
<GID>1099</GID>
<name>clock</name></connection>
<intersection>769.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>769.5,-247.5,825,-247.5</points>
<connection>
<GID>1098</GID>
<name>clock</name></connection>
<intersection>769.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>769.5,-226.5,799,-226.5</points>
<connection>
<GID>1100</GID>
<name>clock</name></connection>
<intersection>769.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>769.5,-210,783,-210</points>
<connection>
<GID>1102</GID>
<name>clock</name></connection>
<intersection>769.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>835.5,-251.5,835.5,-196.5</points>
<connection>
<GID>1114</GID>
<name>OUT_0</name></connection>
<intersection>-251.5 7</intersection>
<intersection>-241.5 10</intersection>
<intersection>-230.5 12</intersection>
<intersection>-221.5 9</intersection>
<intersection>-214 3</intersection>
<intersection>-206.5 8</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>786,-214,835.5,-214</points>
<connection>
<GID>1102</GID>
<name>clear</name></connection>
<intersection>835.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>828,-251.5,835.5,-251.5</points>
<connection>
<GID>1098</GID>
<name>clear</name></connection>
<intersection>835.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>777,-206.5,835.5,-206.5</points>
<connection>
<GID>1103</GID>
<name>clear</name></connection>
<intersection>835.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>794.5,-221.5,835.5,-221.5</points>
<connection>
<GID>1101</GID>
<name>clear</name></connection>
<intersection>835.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>815,-241.5,835.5,-241.5</points>
<connection>
<GID>1099</GID>
<name>clear</name></connection>
<intersection>835.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>802,-230.5,835.5,-230.5</points>
<connection>
<GID>1100</GID>
<name>clear</name></connection>
<intersection>835.5 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-264.58,-1193.57,959.42,-1798.57</PageViewport>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW</type>
<position>273,-524.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>clear</ID>1596 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_OR2</type>
<position>323,-283</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>1410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>193.5,-106</position>
<gparam>LABEL_TEXT Keep Off before setting value and then turn it on</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AE_OR2</type>
<position>324,-567</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>BE_JKFF_LOW_NT</type>
<position>305,-410</position>
<input>
<ID>J</ID>1843 </input>
<output>
<ID>Q</ID>2 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>328,-393.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>293 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND4</type>
<position>473,-252.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>30 </input>
<input>
<ID>IN_3</ID>31 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_OR2</type>
<position>342,-400</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>461 </input>
<output>
<ID>OUT</ID>1842 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>325,-415</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>366,-400</position>
<input>
<ID>N_in0</ID>1844 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AE_DFF_LOW</type>
<position>286.5,-524.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>93 </output>
<input>
<ID>clear</ID>1596 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>15</ID>
<type>BE_JKFF_LOW_NT</type>
<position>194,-717.5</position>
<input>
<ID>J</ID>13 </input>
<output>
<ID>Q</ID>147 </output>
<input>
<ID>clear</ID>13 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>183.5,-727.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>333,-497</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR2</type>
<position>330.5,-746.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>176,-723.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_OR2</type>
<position>338.5,-945.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>348.5,-491.5</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>361,-1167.5</position>
<input>
<ID>N_in0</ID>211 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>201,-719.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR2</type>
<position>334,-1167.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>301.5,-524.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>94 </output>
<input>
<ID>clear</ID>1596 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>349,-483.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_OR2</type>
<position>335.5,-1401.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_DFF_LOW</type>
<position>312,-524.5</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>95 </output>
<input>
<ID>clear</ID>1596 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>325,-524.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>clear</ID>1596 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>358.5,-1401</position>
<input>
<ID>N_in0</ID>222 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>350,-475.5</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>224,-725.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>350.5,-465</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_SMALL_INVERTER</type>
<position>264,-532</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>373.5,-1629</position>
<input>
<ID>N_in0</ID>234 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>BE_JKFF_LOW_NT</type>
<position>212,-926</position>
<input>
<ID>J</ID>149 </input>
<output>
<ID>Q</ID>153 </output>
<input>
<ID>clear</ID>149 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_OR2</type>
<position>344.5,-1628.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>529 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>350,-454</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>201.5,-936</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>BA_NAND2</type>
<position>487.5,-268.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_SMALL_INVERTER</type>
<position>194,-932</position>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>219,-928</position>
<input>
<ID>N_in0</ID>150 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AE_SMALL_INVERTER</type>
<position>279,-532</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AI_XOR2</type>
<position>337,-568</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>242,-934</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>355,-562</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>BE_JKFF_LOW_NT</type>
<position>210.5,-1149</position>
<input>
<ID>J</ID>155 </input>
<output>
<ID>Q</ID>159 </output>
<input>
<ID>clear</ID>155 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_JKFF_LOW_NT</type>
<position>311,-579</position>
<input>
<ID>J</ID>29 </input>
<output>
<ID>Q</ID>79 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_SMALL_INVERTER</type>
<position>294,-532</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_AND2</type>
<position>200,-1159</position>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_SMALL_INVERTER</type>
<position>305.5,-531.5</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>119,-126.5</position>
<output>
<ID>OUT_0</ID>2139 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>167.5,-288.5</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>163,-131</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AE_SMALL_INVERTER</type>
<position>318.5,-532</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_SMALL_INVERTER</type>
<position>331.5,-531.5</position>
<input>
<ID>IN_0</ID>96 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1611</ID>
<type>AI_XOR2</type>
<position>338,-283.5</position>
<input>
<ID>IN_0</ID>1410 </input>
<input>
<ID>IN_1</ID>1411 </input>
<output>
<ID>OUT</ID>1412 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND4</type>
<position>282,-548.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>102 </input>
<input>
<ID>IN_2</ID>100 </input>
<input>
<ID>IN_3</ID>99 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_DFF_LOW</type>
<position>263,-362.5</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clear</ID>1584 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1613</ID>
<type>BA_NAND2</type>
<position>454,-268.5</position>
<input>
<ID>IN_0</ID>1412 </input>
<input>
<ID>IN_1</ID>1411 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_DFF_LOW</type>
<position>276.5,-362.5</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>clear</ID>1584 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>172.5,-418</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-362.5</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clear</ID>1584 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>302,-362.5</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clear</ID>1584 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_DFF_LOW</type>
<position>315,-362.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>72 </output>
<input>
<ID>clear</ID>1584 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND2</type>
<position>318.5,-547.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_SMALL_INVERTER</type>
<position>254,-370</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>296,-570.5</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_SMALL_INVERTER</type>
<position>269,-370</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>284,-370</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>295.5,-369.5</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>308.5,-370</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>290 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_SMALL_INVERTER</type>
<position>321.5,-369.5</position>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>292 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AI_XOR2</type>
<position>253,-515.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AI_XOR2</type>
<position>266.5,-515.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AI_XOR2</type>
<position>279.5,-515.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AI_XOR2</type>
<position>292.5,-515.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AI_XOR2</type>
<position>305,-516</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>330.5,-583</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AI_XOR2</type>
<position>317.5,-516</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>123 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,-1155</position>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>109.5,-396</position>
<gparam>LABEL_TEXT Zone 3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>335.5,-679</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>BE_JKFF_LOW_NT</type>
<position>232,-478.5</position>
<input>
<ID>J</ID>112 </input>
<output>
<ID>Q</ID>113 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>125</ID>
<type>BE_JKFF_LOW_NT</type>
<position>219,-468.5</position>
<input>
<ID>J</ID>114 </input>
<output>
<ID>Q</ID>115 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>126</ID>
<type>BE_JKFF_LOW_NT</type>
<position>206,-457.5</position>
<input>
<ID>J</ID>116 </input>
<output>
<ID>Q</ID>117 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>127</ID>
<type>AI_XOR2</type>
<position>309.5,-563.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>BE_JKFF_LOW_NT</type>
<position>198.5,-448.5</position>
<input>
<ID>J</ID>118 </input>
<output>
<ID>Q</ID>119 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>130</ID>
<type>BE_JKFF_LOW_NT</type>
<position>190,-441</position>
<input>
<ID>J</ID>120 </input>
<output>
<ID>Q</ID>121 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>351,-283</position>
<input>
<ID>N_in0</ID>1412 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>BE_JKFF_LOW_NT</type>
<position>181,-433.5</position>
<input>
<ID>J</ID>122 </input>
<output>
<ID>Q</ID>123 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>137</ID>
<type>CC_PULSE</type>
<position>173,-425.5</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>239.5,-425.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND2</type>
<position>167,-476.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_AND2</type>
<position>166.5,-466.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_AND2</type>
<position>165,-455.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>164.5,-446.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>163.5,-439</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND2</type>
<position>162.5,-431.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_DFF_LOW</type>
<position>257,-524</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>90 </output>
<input>
<ID>clear</ID>1596 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>217.5,-1151</position>
<input>
<ID>N_in0</ID>156 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND2</type>
<position>345.5,-667</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND2</type>
<position>345.5,-658.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>240.5,-1157</position>
<input>
<ID>IN_0</ID>460 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>AI_XOR2</type>
<position>300,-276.5</position>
<input>
<ID>IN_0</ID>325 </input>
<input>
<ID>IN_1</ID>326 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>346.5,-651</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>BE_JKFF_LOW_NT</type>
<position>212.5,-1382.5</position>
<input>
<ID>J</ID>161 </input>
<output>
<ID>Q</ID>165 </output>
<input>
<ID>clear</ID>161 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>347,-642</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>BE_JKFF_LOW_NT</type>
<position>319,-764.5</position>
<input>
<ID>J</ID>145 </input>
<output>
<ID>Q</ID>169 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_AND2</type>
<position>347.5,-634</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND2</type>
<position>202,-1392.5</position>
<input>
<ID>IN_0</ID>512 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>AI_XOR2</type>
<position>345,-747</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_AND2</type>
<position>328.5,-774</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>365.5,-747</position>
<input>
<ID>N_in0</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AE_SMALL_INVERTER</type>
<position>194.5,-1388.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>169</ID>
<type>BA_NAND2</type>
<position>504,-269</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>348,-845.5</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>219.5,-1384.5</position>
<input>
<ID>N_in0</ID>162 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND2</type>
<position>360,-837</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>360,-827</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>242.5,-1390.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>361.5,-820</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>BE_JKFF_LOW_NT</type>
<position>235,-1611</position>
<input>
<ID>J</ID>167 </input>
<output>
<ID>Q</ID>1569 </output>
<input>
<ID>clear</ID>167 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>362,-810.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND2</type>
<position>224.5,-1621</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>1568 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_AND2</type>
<position>362.5,-803.5</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>AE_SMALL_INVERTER</type>
<position>217,-1617</position>
<input>
<ID>IN_0</ID>166 </input>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>AI_XOR2</type>
<position>350,-946</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>GA_LED</type>
<position>242,-1613</position>
<input>
<ID>N_in0</ID>168 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>364,-945.5</position>
<input>
<ID>N_in0</ID>179 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>BA_NAND2</type>
<position>519,-269.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND2</type>
<position>265,-1619</position>
<input>
<ID>IN_0</ID>548 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>1568 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>BE_JKFF_LOW_NT</type>
<position>327,-961</position>
<input>
<ID>J</ID>178 </input>
<output>
<ID>Q</ID>180 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND2</type>
<position>341.5,-969.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND2</type>
<position>339,-1104</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_AND2</type>
<position>350,-1098</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_DFF_LOW</type>
<position>281,-706.5</position>
<input>
<ID>IN_0</ID>185 </input>
<output>
<ID>OUT_0</ID>191 </output>
<input>
<ID>clear</ID>147 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>197</ID>
<type>AE_DFF_LOW</type>
<position>294.5,-706.5</position>
<input>
<ID>IN_0</ID>186 </input>
<output>
<ID>OUT_0</ID>192 </output>
<input>
<ID>clear</ID>147 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>198</ID>
<type>AE_DFF_LOW</type>
<position>309.5,-706.5</position>
<input>
<ID>IN_0</ID>187 </input>
<output>
<ID>OUT_0</ID>193 </output>
<input>
<ID>clear</ID>147 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_DFF_LOW</type>
<position>320,-706.5</position>
<input>
<ID>IN_0</ID>188 </input>
<output>
<ID>OUT_0</ID>194 </output>
<input>
<ID>clear</ID>147 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_DFF_LOW</type>
<position>333,-706.5</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUT_0</ID>195 </output>
<input>
<ID>clear</ID>147 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>201</ID>
<type>AE_SMALL_INVERTER</type>
<position>272,-714</position>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_SMALL_INVERTER</type>
<position>287,-714</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_SMALL_INVERTER</type>
<position>302,-714</position>
<input>
<ID>IN_0</ID>192 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_SMALL_INVERTER</type>
<position>313.5,-713.5</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>AE_SMALL_INVERTER</type>
<position>326.5,-714</position>
<input>
<ID>IN_0</ID>194 </input>
<output>
<ID>OUT_0</ID>200 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>339.5,-713.5</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>201 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_AND4</type>
<position>290,-730.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>198 </input>
<input>
<ID>IN_2</ID>197 </input>
<input>
<ID>IN_3</ID>196 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>180.5,-600</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND2</type>
<position>326.5,-729.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>304,-752.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AI_XOR2</type>
<position>261,-697.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AI_XOR2</type>
<position>274.5,-697.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AI_XOR2</type>
<position>287.5,-697.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>245 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AI_XOR2</type>
<position>300.5,-697.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AI_XOR2</type>
<position>313,-698</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_AND2</type>
<position>350,-1088.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>218</ID>
<type>AI_XOR2</type>
<position>325.5,-698</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>251 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>122,-574</position>
<gparam>LABEL_TEXT Zone 4</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>351,-1079</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>BE_JKFF_LOW_NT</type>
<position>240,-660.5</position>
<input>
<ID>J</ID>232 </input>
<output>
<ID>Q</ID>241 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>223</ID>
<type>BE_JKFF_LOW_NT</type>
<position>227,-650.5</position>
<input>
<ID>J</ID>242 </input>
<output>
<ID>Q</ID>243 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>224</ID>
<type>BE_JKFF_LOW_NT</type>
<position>214,-639.5</position>
<input>
<ID>J</ID>244 </input>
<output>
<ID>Q</ID>245 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>225</ID>
<type>AI_XOR2</type>
<position>317.5,-745.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>BE_JKFF_LOW_NT</type>
<position>206.5,-630.5</position>
<input>
<ID>J</ID>246 </input>
<output>
<ID>Q</ID>247 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>227</ID>
<type>BE_JKFF_LOW_NT</type>
<position>198,-623</position>
<input>
<ID>J</ID>248 </input>
<output>
<ID>Q</ID>249 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>228</ID>
<type>BE_JKFF_LOW_NT</type>
<position>189,-615.5</position>
<input>
<ID>J</ID>250 </input>
<output>
<ID>Q</ID>251 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>229</ID>
<type>CC_PULSE</type>
<position>180.5,-607.5</position>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>175,-658.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_AND2</type>
<position>174.5,-648.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>173,-637.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_AND2</type>
<position>172.5,-628.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>246 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>351.5,-1070.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_AND2</type>
<position>352.5,-1062</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AI_XOR2</type>
<position>346.5,-1168.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AI_XOR2</type>
<position>-241,173</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>1572 </input>
<output>
<ID>OUT</ID>1576 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>BE_JKFF_LOW_NT</type>
<position>321.5,-1186</position>
<input>
<ID>J</ID>210 </input>
<output>
<ID>Q</ID>212 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_AND2</type>
<position>335.5,-1187.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1783</ID>
<type>BE_JKFF_LOW_NT</type>
<position>222,-254.5</position>
<input>
<ID>J</ID>1574 </input>
<output>
<ID>Q</ID>1571 </output>
<input>
<ID>clear</ID>1574 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>1575 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_AND2</type>
<position>339.5,-1343.5</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1785</ID>
<type>AA_AND2</type>
<position>161.5,-271</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>1578 </input>
<output>
<ID>OUT</ID>1573 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_AND2</type>
<position>350.5,-1334</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>171.5,-621</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_AND2</type>
<position>350,-1324.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>1570 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1789</ID>
<type>AE_SMALL_INVERTER</type>
<position>204,-260.5</position>
<input>
<ID>IN_0</ID>1573 </input>
<output>
<ID>OUT_0</ID>1574 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>350.5,-1316</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1791</ID>
<type>GA_LED</type>
<position>229,-256.5</position>
<input>
<ID>N_in0</ID>1575 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>AA_AND2</type>
<position>350.5,-1307.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1793</ID>
<type>AA_TOGGLE</type>
<position>196,-111</position>
<output>
<ID>OUT_0</ID>1577 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_AND2</type>
<position>351,-1300</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1795</ID>
<type>AA_AND2</type>
<position>172.5,-267</position>
<input>
<ID>IN_0</ID>325 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>1578 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1796</ID>
<type>BE_JKFF_LOW_NT</type>
<position>219,-379</position>
<input>
<ID>J</ID>1580 </input>
<output>
<ID>Q</ID>1584 </output>
<input>
<ID>clear</ID>1580 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>1581 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1797</ID>
<type>AA_AND2</type>
<position>149,-390</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>1583 </input>
<output>
<ID>OUT</ID>1579 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1798</ID>
<type>AE_SMALL_INVERTER</type>
<position>142,-388</position>
<input>
<ID>IN_0</ID>1579 </input>
<output>
<ID>OUT_0</ID>1580 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>261</ID>
<type>BA_NAND2</type>
<position>533,-269.5</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1799</ID>
<type>GA_LED</type>
<position>226,-381</position>
<input>
<ID>N_in0</ID>1581 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AI_XOR2</type>
<position>348,-1401.5</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1801</ID>
<type>AA_AND2</type>
<position>161,-389</position>
<input>
<ID>IN_0</ID>293 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>1583 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>BA_NAND2</type>
<position>546,-269.5</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>BE_JKFF_LOW_NT</type>
<position>326,-1420.5</position>
<input>
<ID>J</ID>221 </input>
<output>
<ID>Q</ID>223 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_AND2</type>
<position>341.5,-1425</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>529 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1808</ID>
<type>BE_JKFF_LOW_NT</type>
<position>195,-550</position>
<input>
<ID>J</ID>1592 </input>
<output>
<ID>Q</ID>1596 </output>
<input>
<ID>clear</ID>1592 </input>
<input>
<ID>clock</ID>397 </input>
<output>
<ID>nQ</ID>1593 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND2</type>
<position>357,-1565</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1809</ID>
<type>AA_AND2</type>
<position>184.5,-560</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>1595 </input>
<output>
<ID>OUT</ID>1591 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1810</ID>
<type>AE_SMALL_INVERTER</type>
<position>177,-556</position>
<input>
<ID>IN_0</ID>1591 </input>
<output>
<ID>OUT_0</ID>1592 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_AND2</type>
<position>369,-1556.5</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1811</ID>
<type>GA_LED</type>
<position>202,-552</position>
<input>
<ID>N_in0</ID>1593 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>AA_AND2</type>
<position>370.5,-1546.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1813</ID>
<type>AA_AND2</type>
<position>225,-558</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>1577 </input>
<output>
<ID>OUT</ID>1595 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1814</ID>
<type>AA_TOGGLE</type>
<position>131,-126</position>
<output>
<ID>OUT_0</ID>2140 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_AND2</type>
<position>170.5,-613.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1816</ID>
<type>AA_LABEL</type>
<position>134.5,-121</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>AE_DFF_LOW</type>
<position>265,-706</position>
<input>
<ID>IN_0</ID>184 </input>
<output>
<ID>OUT_0</ID>190 </output>
<input>
<ID>clear</ID>147 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>279</ID>
<type>AE_DFF_LOW</type>
<position>291.5,-905.5</position>
<input>
<ID>IN_0</ID>257 </input>
<output>
<ID>OUT_0</ID>263 </output>
<input>
<ID>clear</ID>153 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1818</ID>
<type>AI_XOR2</type>
<position>123.5,-136</position>
<input>
<ID>IN_0</ID>2140 </input>
<input>
<ID>IN_1</ID>2139 </input>
<output>
<ID>OUT</ID>304 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AE_DFF_LOW</type>
<position>305,-905.5</position>
<input>
<ID>IN_0</ID>258 </input>
<output>
<ID>OUT_0</ID>264 </output>
<input>
<ID>clear</ID>153 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>281</ID>
<type>AE_DFF_LOW</type>
<position>320,-905.5</position>
<input>
<ID>IN_0</ID>259 </input>
<output>
<ID>OUT_0</ID>265 </output>
<input>
<ID>clear</ID>153 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1820</ID>
<type>AI_XOR2</type>
<position>128.5,-288</position>
<input>
<ID>IN_0</ID>2142 </input>
<input>
<ID>IN_1</ID>2141 </input>
<output>
<ID>OUT</ID>461 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AE_DFF_LOW</type>
<position>330.5,-905.5</position>
<input>
<ID>IN_0</ID>260 </input>
<output>
<ID>OUT_0</ID>266 </output>
<input>
<ID>clear</ID>153 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>283</ID>
<type>AE_DFF_LOW</type>
<position>343.5,-905.5</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>267 </output>
<input>
<ID>clear</ID>153 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1822</ID>
<type>AA_TOGGLE</type>
<position>130,-279.5</position>
<output>
<ID>OUT_0</ID>2142 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>284</ID>
<type>AE_SMALL_INVERTER</type>
<position>282.5,-913</position>
<input>
<ID>IN_0</ID>262 </input>
<output>
<ID>OUT_0</ID>268 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>285</ID>
<type>AE_SMALL_INVERTER</type>
<position>297.5,-913</position>
<input>
<ID>IN_0</ID>263 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1824</ID>
<type>AA_LABEL</type>
<position>131,-275.5</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>AE_SMALL_INVERTER</type>
<position>312.5,-913</position>
<input>
<ID>IN_0</ID>264 </input>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1825</ID>
<type>AI_XOR2</type>
<position>119.5,-411.5</position>
<input>
<ID>IN_0</ID>2144 </input>
<input>
<ID>IN_1</ID>2143 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>AE_SMALL_INVERTER</type>
<position>324,-912.5</position>
<input>
<ID>IN_0</ID>265 </input>
<output>
<ID>OUT_0</ID>271 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1826</ID>
<type>AA_TOGGLE</type>
<position>121,-403</position>
<output>
<ID>OUT_0</ID>2144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_SMALL_INVERTER</type>
<position>337,-913</position>
<input>
<ID>IN_0</ID>266 </input>
<output>
<ID>OUT_0</ID>272 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1827</ID>
<type>AA_LABEL</type>
<position>122,-399</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>350,-912.5</position>
<input>
<ID>IN_0</ID>267 </input>
<output>
<ID>OUT_0</ID>273 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1828</ID>
<type>AA_TOGGLE</type>
<position>114.5,-403</position>
<output>
<ID>OUT_0</ID>2143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1829</ID>
<type>AI_XOR2</type>
<position>133,-588</position>
<input>
<ID>IN_0</ID>2146 </input>
<input>
<ID>IN_1</ID>2145 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_AND4</type>
<position>300.5,-929.5</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>270 </input>
<input>
<ID>IN_2</ID>269 </input>
<input>
<ID>IN_3</ID>268 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1830</ID>
<type>AA_TOGGLE</type>
<position>136,-579</position>
<output>
<ID>OUT_0</ID>2146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>191,-799</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1831</ID>
<type>AA_LABEL</type>
<position>142,-575</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_AND2</type>
<position>337,-928.5</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1832</ID>
<type>AA_TOGGLE</type>
<position>129,-579</position>
<output>
<ID>OUT_0</ID>2145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_AND2</type>
<position>314.5,-951.5</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1833</ID>
<type>AI_XOR2</type>
<position>152.5,-785</position>
<input>
<ID>IN_0</ID>2148 </input>
<input>
<ID>IN_1</ID>2147 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>AI_XOR2</type>
<position>271.5,-896.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>278 </input>
<output>
<ID>OUT</ID>256 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1834</ID>
<type>AA_TOGGLE</type>
<position>154,-776.5</position>
<output>
<ID>OUT_0</ID>2148 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>296</ID>
<type>AI_XOR2</type>
<position>285,-896.5</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>280 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1835</ID>
<type>AA_LABEL</type>
<position>155,-772.5</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>AI_XOR2</type>
<position>298,-896.5</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>282 </input>
<output>
<ID>OUT</ID>258 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1836</ID>
<type>AA_TOGGLE</type>
<position>147.5,-776.5</position>
<output>
<ID>OUT_0</ID>2147 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>298</ID>
<type>AI_XOR2</type>
<position>311,-896.5</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1837</ID>
<type>AI_XOR2</type>
<position>146,-1002.5</position>
<input>
<ID>IN_0</ID>2150 </input>
<input>
<ID>IN_1</ID>2149 </input>
<output>
<ID>OUT</ID>296 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>AI_XOR2</type>
<position>323.5,-897</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>286 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1838</ID>
<type>AA_TOGGLE</type>
<position>147.5,-994</position>
<output>
<ID>OUT_0</ID>2150 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND2</type>
<position>371,-1537</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1839</ID>
<type>AA_LABEL</type>
<position>148.5,-990</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>AI_XOR2</type>
<position>336,-897</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1840</ID>
<type>AA_TOGGLE</type>
<position>141,-994</position>
<output>
<ID>OUT_0</ID>2149 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1841</ID>
<type>AI_XOR2</type>
<position>147,-1244.5</position>
<input>
<ID>IN_0</ID>2152 </input>
<input>
<ID>IN_1</ID>2151 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>140.5,-768.5</position>
<gparam>LABEL_TEXT Zone 5</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1842</ID>
<type>AA_TOGGLE</type>
<position>148.5,-1236</position>
<output>
<ID>OUT_0</ID>2152 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>370.5,-1528.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1843</ID>
<type>AA_LABEL</type>
<position>149.5,-1232</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>BE_JKFF_LOW_NT</type>
<position>250.5,-859.5</position>
<input>
<ID>J</ID>277 </input>
<output>
<ID>Q</ID>278 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1844</ID>
<type>AA_TOGGLE</type>
<position>142,-1236</position>
<output>
<ID>OUT_0</ID>2151 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>306</ID>
<type>BE_JKFF_LOW_NT</type>
<position>237.5,-849.5</position>
<input>
<ID>J</ID>279 </input>
<output>
<ID>Q</ID>280 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1845</ID>
<type>AI_XOR2</type>
<position>154,-1458</position>
<input>
<ID>IN_0</ID>2154 </input>
<input>
<ID>IN_1</ID>2153 </input>
<output>
<ID>OUT</ID>529 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>BE_JKFF_LOW_NT</type>
<position>224.5,-838.5</position>
<input>
<ID>J</ID>281 </input>
<output>
<ID>Q</ID>282 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1846</ID>
<type>AA_TOGGLE</type>
<position>155.5,-1449.5</position>
<output>
<ID>OUT_0</ID>2154 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>308</ID>
<type>AI_XOR2</type>
<position>328,-944.5</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1847</ID>
<type>AA_LABEL</type>
<position>156.5,-1445.5</position>
<gparam>LABEL_TEXT Disable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>BE_JKFF_LOW_NT</type>
<position>217,-829.5</position>
<input>
<ID>J</ID>283 </input>
<output>
<ID>Q</ID>284 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1848</ID>
<type>AA_TOGGLE</type>
<position>149,-1449.5</position>
<output>
<ID>OUT_0</ID>2153 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>310</ID>
<type>BE_JKFF_LOW_NT</type>
<position>208.5,-822</position>
<input>
<ID>J</ID>285 </input>
<output>
<ID>Q</ID>286 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>311</ID>
<type>BE_JKFF_LOW_NT</type>
<position>199.5,-814.5</position>
<input>
<ID>J</ID>287 </input>
<output>
<ID>Q</ID>288 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1850</ID>
<type>GA_LED</type>
<position>154,-126</position>
<input>
<ID>N_in0</ID>2140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>CC_PULSE</type>
<position>191.5,-806.5</position>
<output>
<ID>OUT_0</ID>289 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>185.5,-857.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1853</ID>
<type>GA_LED</type>
<position>142,-280.5</position>
<input>
<ID>N_in0</ID>2142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AA_AND2</type>
<position>185,-847.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1854</ID>
<type>GA_LED</type>
<position>132.5,-403.5</position>
<input>
<ID>N_in0</ID>2144 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>183.5,-836.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1855</ID>
<type>GA_LED</type>
<position>148.5,-581</position>
<input>
<ID>N_in0</ID>2146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>AA_AND2</type>
<position>183,-827.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1856</ID>
<type>GA_LED</type>
<position>165.5,-779</position>
<input>
<ID>N_in0</ID>2148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AA_AND2</type>
<position>182,-820</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>285 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1857</ID>
<type>GA_LED</type>
<position>158,-997.5</position>
<input>
<ID>N_in0</ID>2150 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>181,-812.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1858</ID>
<type>GA_LED</type>
<position>159.5,-1238.5</position>
<input>
<ID>N_in0</ID>2152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AE_DFF_LOW</type>
<position>275.5,-905</position>
<input>
<ID>IN_0</ID>256 </input>
<output>
<ID>OUT_0</ID>262 </output>
<input>
<ID>clear</ID>153 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1859</ID>
<type>GA_LED</type>
<position>165.5,-1452.5</position>
<input>
<ID>N_in0</ID>2154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>321</ID>
<type>AE_DFF_LOW</type>
<position>285,-1127.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>327 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_DFF_LOW</type>
<position>299,-1127.5</position>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>328 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_DFF_LOW</type>
<position>313.5,-1127.5</position>
<input>
<ID>IN_0</ID>302 </input>
<output>
<ID>OUT_0</ID>329 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_DFF_LOW</type>
<position>324,-1127.5</position>
<input>
<ID>IN_0</ID>303 </input>
<output>
<ID>OUT_0</ID>400 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_AND4</type>
<position>272,-386.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>77 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>326</ID>
<type>AA_AND2</type>
<position>308.5,-385.5</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>290 </input>
<output>
<ID>OUT</ID>294 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>287.5,-403.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>293 </input>
<output>
<ID>OUT</ID>1843 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>AI_XOR2</type>
<position>243,-353.5</position>
<input>
<ID>IN_0</ID>1836 </input>
<input>
<ID>IN_1</ID>594 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AI_XOR2</type>
<position>256.5,-353.5</position>
<input>
<ID>IN_0</ID>1837 </input>
<input>
<ID>IN_1</ID>596 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AI_XOR2</type>
<position>269.5,-353.5</position>
<input>
<ID>IN_0</ID>1838 </input>
<input>
<ID>IN_1</ID>598 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AI_XOR2</type>
<position>282.5,-353.5</position>
<input>
<ID>IN_0</ID>1839 </input>
<input>
<ID>IN_1</ID>600 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AI_XOR2</type>
<position>295,-354</position>
<input>
<ID>IN_0</ID>1840 </input>
<input>
<ID>IN_1</ID>602 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AI_XOR2</type>
<position>307.5,-354</position>
<input>
<ID>IN_0</ID>1841 </input>
<input>
<ID>IN_1</ID>604 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>334</ID>
<type>AE_DFF_LOW</type>
<position>247,-362</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clear</ID>1584 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_DFF_LOW</type>
<position>337,-1127.5</position>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>407 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_SMALL_INVERTER</type>
<position>276,-1135</position>
<input>
<ID>IN_0</ID>306 </input>
<output>
<ID>OUT_0</ID>408 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_AND2</type>
<position>157.5,-189.5</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>470 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_SMALL_INVERTER</type>
<position>291,-1135</position>
<input>
<ID>IN_0</ID>327 </input>
<output>
<ID>OUT_0</ID>455 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>339</ID>
<type>AE_SMALL_INVERTER</type>
<position>306,-1135</position>
<input>
<ID>IN_0</ID>328 </input>
<output>
<ID>OUT_0</ID>456 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>157,-179.5</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AA_AND2</type>
<position>155.5,-168.5</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>474 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>AE_SMALL_INVERTER</type>
<position>317.5,-1134.5</position>
<input>
<ID>IN_0</ID>329 </input>
<output>
<ID>OUT_0</ID>457 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_AND2</type>
<position>155,-159.5</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>476 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_SMALL_INVERTER</type>
<position>330.5,-1135</position>
<input>
<ID>IN_0</ID>400 </input>
<output>
<ID>OUT_0</ID>458 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>345</ID>
<type>AE_SMALL_INVERTER</type>
<position>343.5,-1134.5</position>
<input>
<ID>IN_0</ID>407 </input>
<output>
<ID>OUT_0</ID>459 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>346</ID>
<type>AA_AND2</type>
<position>154,-152</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>478 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>AA_AND2</type>
<position>153,-144.5</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>480 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>-133.5,-147.5</position>
<gparam>LABEL_TEXT Checking condition for 60</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>AA_TOGGLE</type>
<position>-264,-8.5</position>
<output>
<ID>OUT_0</ID>331 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_LABEL</type>
<position>68,-66.5</position>
<gparam>LABEL_TEXT Problematic Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>BA_NAND4</type>
<position>45,-11.5</position>
<input>
<ID>IN_0</ID>348 </input>
<input>
<ID>IN_1</ID>352 </input>
<input>
<ID>IN_2</ID>356 </input>
<input>
<ID>IN_3</ID>361 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_DFF_LOW</type>
<position>-154,-81.5</position>
<input>
<ID>IN_0</ID>339 </input>
<output>
<ID>OUT_0</ID>344 </output>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>355</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-172,-37</position>
<input>
<ID>J</ID>367 </input>
<input>
<ID>K</ID>369 </input>
<output>
<ID>Q</ID>339 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>360 </input>
<output>
<ID>nQ</ID>340 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>357</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-122.5,-37.5</position>
<input>
<ID>J</ID>379 </input>
<input>
<ID>K</ID>380 </input>
<output>
<ID>Q</ID>343 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>360 </input>
<output>
<ID>nQ</ID>346 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>358</ID>
<type>AE_DFF_LOW</type>
<position>-111,-81</position>
<input>
<ID>IN_0</ID>343 </input>
<output>
<ID>OUT_0</ID>362 </output>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>359</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-96.5,-37</position>
<input>
<ID>J</ID>381 </input>
<input>
<ID>K</ID>382 </input>
<output>
<ID>Q</ID>348 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>360 </input>
<output>
<ID>nQ</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>361</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-66.5,-37.5</position>
<input>
<ID>J</ID>383 </input>
<input>
<ID>K</ID>384 </input>
<output>
<ID>Q</ID>352 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>360 </input>
<output>
<ID>nQ</ID>353 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>363</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-28,-39.5</position>
<input>
<ID>J</ID>385 </input>
<input>
<ID>K</ID>386 </input>
<output>
<ID>Q</ID>356 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>360 </input>
<output>
<ID>nQ</ID>357 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>365</ID>
<type>BE_JKFF_LOW_NT</type>
<position>20.5,-40</position>
<input>
<ID>J</ID>387 </input>
<input>
<ID>K</ID>388 </input>
<output>
<ID>Q</ID>361 </output>
<input>
<ID>clear</ID>338 </input>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_DFF_LOW</type>
<position>-81.5,-81</position>
<input>
<ID>IN_0</ID>348 </input>
<output>
<ID>OUT_0</ID>363 </output>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_AND2</type>
<position>-155.5,-28</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>339 </input>
<output>
<ID>OUT</ID>341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_DFF_LOW</type>
<position>247.5,-237</position>
<input>
<ID>IN_0</ID>307 </input>
<output>
<ID>OUT_0</ID>313 </output>
<input>
<ID>clear</ID>1571 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_AND2</type>
<position>-156.5,-45.5</position>
<input>
<ID>IN_0</ID>340 </input>
<input>
<ID>IN_1</ID>396 </input>
<output>
<ID>OUT</ID>342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_AND2</type>
<position>-114.5,-28</position>
<input>
<ID>IN_0</ID>341 </input>
<input>
<ID>IN_1</ID>343 </input>
<output>
<ID>OUT</ID>345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_AND2</type>
<position>-112,-46.5</position>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>342 </input>
<output>
<ID>OUT</ID>347 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>-85,-29.5</position>
<input>
<ID>IN_0</ID>345 </input>
<input>
<ID>IN_1</ID>348 </input>
<output>
<ID>OUT</ID>349 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_AND2</type>
<position>-82.5,-48</position>
<input>
<ID>IN_0</ID>351 </input>
<input>
<ID>IN_1</ID>347 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_AND2</type>
<position>-58.5,-30.5</position>
<input>
<ID>IN_0</ID>349 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_AND2</type>
<position>-57,-48</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>350 </input>
<output>
<ID>OUT</ID>355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>AA_AND2</type>
<position>-11.5,-29.5</position>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>356 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND2</type>
<position>-11,-47</position>
<input>
<ID>IN_0</ID>357 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>359 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AE_DFF_LOW</type>
<position>-53,-81</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>364 </output>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_OR2</type>
<position>-141.5,-37.5</position>
<input>
<ID>IN_0</ID>341 </input>
<input>
<ID>IN_1</ID>342 </input>
<output>
<ID>OUT</ID>379 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AE_DFF_LOW</type>
<position>-7,-81</position>
<input>
<ID>IN_0</ID>356 </input>
<output>
<ID>OUT_0</ID>365 </output>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>382</ID>
<type>AE_OR2</type>
<position>-105,-36.5</position>
<input>
<ID>IN_0</ID>345 </input>
<input>
<ID>IN_1</ID>347 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_OR2</type>
<position>-76.5,-37</position>
<input>
<ID>IN_0</ID>349 </input>
<input>
<ID>IN_1</ID>350 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>AE_OR2</type>
<position>-47.5,-37.5</position>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>385 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>AE_OR2</type>
<position>-3.5,-38</position>
<input>
<ID>IN_0</ID>358 </input>
<input>
<ID>IN_1</ID>359 </input>
<output>
<ID>OUT</ID>387 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>386</ID>
<type>AE_DFF_LOW</type>
<position>41,-81.5</position>
<input>
<ID>IN_0</ID>361 </input>
<output>
<ID>OUT_0</ID>366 </output>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>387</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>45,-61</position>
<input>
<ID>IN_0</ID>339 </input>
<input>
<ID>IN_1</ID>343 </input>
<input>
<ID>IN_2</ID>348 </input>
<input>
<ID>IN_3</ID>352 </input>
<input>
<ID>IN_4</ID>356 </input>
<input>
<ID>IN_5</ID>361 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>388</ID>
<type>AE_DFF_LOW</type>
<position>-235.5,-45.5</position>
<input>
<ID>IN_0</ID>394 </input>
<output>
<ID>OUTINV_0</ID>396 </output>
<output>
<ID>OUT_0</ID>395 </output>
<input>
<ID>clear</ID>337 </input>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>389</ID>
<type>CC_PULSE</type>
<position>-283,-40</position>
<output>
<ID>OUT_0</ID>392 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>64.5,-91.5</position>
<input>
<ID>IN_0</ID>344 </input>
<input>
<ID>IN_1</ID>362 </input>
<input>
<ID>IN_2</ID>363 </input>
<input>
<ID>IN_3</ID>364 </input>
<input>
<ID>IN_4</ID>365 </input>
<input>
<ID>IN_5</ID>366 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>391</ID>
<type>CC_PULSE</type>
<position>-281.5,-58</position>
<output>
<ID>OUT_0</ID>391 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>392</ID>
<type>EE_VDD</type>
<position>-231,-5</position>
<output>
<ID>OUT_0</ID>390 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>393</ID>
<type>AE_OR2</type>
<position>-244.5,-57</position>
<input>
<ID>IN_0</ID>392 </input>
<input>
<ID>IN_1</ID>391 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>AE_DFF_LOW</type>
<position>263.5,-237.5</position>
<input>
<ID>IN_0</ID>308 </input>
<output>
<ID>OUT_0</ID>314 </output>
<input>
<ID>clear</ID>1571 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>395</ID>
<type>AE_SMALL_INVERTER</type>
<position>-262,-40.5</position>
<input>
<ID>IN_0</ID>392 </input>
<output>
<ID>OUT_0</ID>393 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_AND2</type>
<position>-138,-132</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>372 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>397</ID>
<type>AI_XOR2</type>
<position>-247.5,-44.5</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>393 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_LABEL</type>
<position>-277.5,-34</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>399</ID>
<type>AA_AND2</type>
<position>-64,-118.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>374 </input>
<output>
<ID>OUT</ID>375 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>-278.5,-63</position>
<gparam>LABEL_TEXT Decrement</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>AA_AND2</type>
<position>-1,-117</position>
<input>
<ID>IN_0</ID>376 </input>
<input>
<ID>IN_1</ID>377 </input>
<output>
<ID>OUT</ID>378 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>AI_XOR2</type>
<position>-187.5,-26</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>369 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>AE_DFF_LOW</type>
<position>277,-237.5</position>
<input>
<ID>IN_0</ID>309 </input>
<output>
<ID>OUT_0</ID>315 </output>
<input>
<ID>clear</ID>1571 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>404</ID>
<type>AI_XOR2</type>
<position>-136.5,-23.5</position>
<input>
<ID>IN_0</ID>379 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>AI_XOR2</type>
<position>-100,-23</position>
<input>
<ID>IN_0</ID>382 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>381 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AI_XOR2</type>
<position>-71.5,-23.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>384 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AI_XOR2</type>
<position>-41.5,-23.5</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AI_XOR2</type>
<position>6,-21.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>388 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND4</type>
<position>-159.5,-154</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>375 </input>
<input>
<ID>IN_2</ID>372 </input>
<input>
<ID>IN_3</ID>396 </input>
<output>
<ID>OUT</ID>368 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_DFF_LOW</type>
<position>292,-237.5</position>
<input>
<ID>IN_0</ID>310 </input>
<output>
<ID>OUT_0</ID>316 </output>
<input>
<ID>clear</ID>1571 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_INVERTER</type>
<position>-144,-109</position>
<input>
<ID>IN_0</ID>339 </input>
<output>
<ID>OUT_0</ID>370 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_INVERTER</type>
<position>-131.5,-110</position>
<input>
<ID>IN_0</ID>343 </input>
<output>
<ID>OUT_0</ID>371 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>413</ID>
<type>AA_INVERTER</type>
<position>-67.5,-109</position>
<input>
<ID>IN_0</ID>348 </input>
<output>
<ID>OUT_0</ID>374 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>414</ID>
<type>AA_INVERTER</type>
<position>-60.5,-109</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>373 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>415</ID>
<type>AE_DFF_LOW</type>
<position>302.5,-237.5</position>
<input>
<ID>IN_0</ID>311 </input>
<output>
<ID>OUT_0</ID>317 </output>
<input>
<ID>clear</ID>1571 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_INVERTER</type>
<position>-3,-108.5</position>
<input>
<ID>IN_0</ID>356 </input>
<output>
<ID>OUT_0</ID>377 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>417</ID>
<type>AA_INVERTER</type>
<position>2.5,-108</position>
<input>
<ID>IN_0</ID>361 </input>
<output>
<ID>OUT_0</ID>376 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>64.5,-101.5</position>
<gparam>LABEL_TEXT Actual Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>419</ID>
<type>AA_AND4</type>
<position>294,-1151.5</position>
<input>
<ID>IN_0</ID>457 </input>
<input>
<ID>IN_1</ID>456 </input>
<input>
<ID>IN_2</ID>455 </input>
<input>
<ID>IN_3</ID>408 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_AND2</type>
<position>-238,-11.5</position>
<input>
<ID>IN_0</ID>390 </input>
<input>
<ID>IN_1</ID>389 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>AA_LABEL</type>
<position>-109,-2</position>
<gparam>LABEL_TEXT Setting Mode</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>AE_DFF_LOW</type>
<position>315.5,-237.5</position>
<input>
<ID>IN_0</ID>312 </input>
<output>
<ID>OUT_0</ID>318 </output>
<input>
<ID>clear</ID>1571 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>-244,1.5</position>
<gparam>LABEL_TEXT On/Off- Settings/Cycle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>AA_LABEL</type>
<position>184.5,-1021</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>AA_LABEL</type>
<position>-271,183</position>
<gparam>LABEL_TEXT Water Button</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>AE_SMALL_INVERTER</type>
<position>254.5,-245</position>
<input>
<ID>IN_0</ID>313 </input>
<output>
<ID>OUT_0</ID>319 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>428</ID>
<type>AA_LABEL</type>
<position>-107,149</position>
<gparam>LABEL_TEXT Buffer Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>AA_LABEL</type>
<position>-165,200.5</position>
<gparam>LABEL_TEXT Seconds Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>430</ID>
<type>AE_SMALL_INVERTER</type>
<position>269.5,-245</position>
<input>
<ID>IN_0</ID>314 </input>
<output>
<ID>OUT_0</ID>320 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>431</ID>
<type>BE_JKFF_LOW_NT</type>
<position>22,87.5</position>
<input>
<ID>J</ID>453 </input>
<input>
<ID>K</ID>1414 </input>
<output>
<ID>Q</ID>398 </output>
<input>
<ID>clear</ID>254 </input>
<input>
<ID>clock</ID>425 </input>
<output>
<ID>nQ</ID>404 </output>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>432</ID>
<type>AA_LABEL</type>
<position>-108.5,127.5</position>
<gparam>LABEL_TEXT Actual Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AE_SMALL_INVERTER</type>
<position>284.5,-245</position>
<input>
<ID>IN_0</ID>315 </input>
<output>
<ID>OUT_0</ID>321 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>-34.5,109</position>
<gparam>LABEL_TEXT Minutes Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AE_SMALL_INVERTER</type>
<position>296,-244.5</position>
<input>
<ID>IN_0</ID>316 </input>
<output>
<ID>OUT_0</ID>322 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>436</ID>
<type>AA_LABEL</type>
<position>28.5,73.5</position>
<gparam>LABEL_TEXT Buffer Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AE_SMALL_INVERTER</type>
<position>309,-245</position>
<input>
<ID>IN_0</ID>317 </input>
<output>
<ID>OUT_0</ID>323 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>438</ID>
<type>AI_XOR2</type>
<position>-92.5,173.5</position>
<input>
<ID>IN_0</ID>404 </input>
<input>
<ID>IN_1</ID>406 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>-88,183.5</position>
<gparam>LABEL_TEXT Both on seconds counter stop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AE_SMALL_INVERTER</type>
<position>322,-244.5</position>
<input>
<ID>IN_0</ID>318 </input>
<output>
<ID>OUT_0</ID>324 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>441</ID>
<type>AA_LABEL</type>
<position>38,44.5</position>
<gparam>LABEL_TEXT Actual Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>AI_XOR2</type>
<position>6.5,85.5</position>
<input>
<ID>IN_0</ID>416 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>AA_INVERTER</type>
<position>15.5,102.5</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>1414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>444</ID>
<type>AA_AND2</type>
<position>-231,150</position>
<input>
<ID>IN_0</ID>453 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>425 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_LABEL</type>
<position>-242,76</position>
<gparam>LABEL_TEXT Abort</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>446</ID>
<type>AE_OR2</type>
<position>-177.5,94</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>402 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>447</ID>
<type>AA_TOGGLE</type>
<position>-244,79.5</position>
<output>
<ID>OUT_0</ID>416 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>448</ID>
<type>AE_OR4</type>
<position>-209.5,102.5</position>
<input>
<ID>IN_0</ID>434 </input>
<input>
<ID>IN_1</ID>433 </input>
<input>
<ID>IN_2</ID>432 </input>
<input>
<ID>IN_3</ID>431 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>449</ID>
<type>AE_OR2</type>
<position>-223.5,97</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>399 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>450</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-218.5,162.5</position>
<input>
<ID>J</ID>453 </input>
<input>
<ID>K</ID>453 </input>
<output>
<ID>Q</ID>424 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>451</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-205,162.5</position>
<input>
<ID>J</ID>424 </input>
<input>
<ID>K</ID>424 </input>
<output>
<ID>Q</ID>426 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>452</ID>
<type>AA_AND2</type>
<position>-230,106.5</position>
<input>
<ID>IN_0</ID>401 </input>
<input>
<ID>IN_1</ID>453 </input>
<output>
<ID>OUT</ID>403 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>453</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-189,162.5</position>
<input>
<ID>J</ID>420 </input>
<input>
<ID>K</ID>420 </input>
<output>
<ID>Q</ID>428 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>454</ID>
<type>AE_OR2</type>
<position>-248.5,109.5</position>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>403 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>455</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-173,162</position>
<input>
<ID>J</ID>421 </input>
<input>
<ID>K</ID>421 </input>
<output>
<ID>Q</ID>427 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>456</ID>
<type>AA_AND4</type>
<position>272.5,-261.5</position>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>321 </input>
<input>
<ID>IN_2</ID>320 </input>
<input>
<ID>IN_3</ID>319 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>457</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-157,161.5</position>
<input>
<ID>J</ID>422 </input>
<input>
<ID>K</ID>422 </input>
<output>
<ID>Q</ID>429 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>458</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-140,161.5</position>
<input>
<ID>J</ID>423 </input>
<input>
<ID>K</ID>423 </input>
<output>
<ID>Q</ID>430 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>459</ID>
<type>AI_XOR2</type>
<position>-107.5,164.5</position>
<input>
<ID>IN_0</ID>416 </input>
<input>
<ID>IN_1</ID>413 </input>
<output>
<ID>OUT</ID>405 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AA_TOGGLE</type>
<position>-255.5,173</position>
<output>
<ID>OUT_0</ID>1572 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>461</ID>
<type>AA_LABEL</type>
<position>-262,116.5</position>
<gparam>LABEL_TEXT Water On/Off</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>462</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-90,89.5</position>
<input>
<ID>J</ID>453 </input>
<input>
<ID>K</ID>453 </input>
<output>
<ID>Q</ID>441 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_AND2</type>
<position>-241,98</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>453 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-76.5,89.5</position>
<input>
<ID>J</ID>441 </input>
<input>
<ID>K</ID>441 </input>
<output>
<ID>Q</ID>442 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>465</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-122.5,148</position>
<input>
<ID>IN_0</ID>424 </input>
<input>
<ID>IN_1</ID>426 </input>
<input>
<ID>IN_2</ID>428 </input>
<input>
<ID>IN_3</ID>427 </input>
<input>
<ID>IN_4</ID>429 </input>
<input>
<ID>IN_5</ID>430 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>466</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-60.5,89.5</position>
<input>
<ID>J</ID>437 </input>
<input>
<ID>K</ID>437 </input>
<output>
<ID>Q</ID>444 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>467</ID>
<type>AA_AND2</type>
<position>309,-260.5</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>468</ID>
<type>GA_LED</type>
<position>-260.5,109.5</position>
<input>
<ID>N_in1</ID>411 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>469</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-44.5,89</position>
<input>
<ID>J</ID>438 </input>
<input>
<ID>K</ID>438 </input>
<output>
<ID>Q</ID>443 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_AND2</type>
<position>286.5,-283.5</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>1411 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>AA_LABEL</type>
<position>-210,91.5</position>
<gparam>LABEL_TEXT Output of Flip-flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>472</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-28.5,89.5</position>
<input>
<ID>J</ID>439 </input>
<input>
<ID>K</ID>439 </input>
<output>
<ID>Q</ID>445 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>473</ID>
<type>BB_CLOCK</type>
<position>-245.5,149</position>
<output>
<ID>CLK</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 3</lparam></gate>
<gate>
<ID>474</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-11.5,89.5</position>
<input>
<ID>J</ID>440 </input>
<input>
<ID>K</ID>440 </input>
<output>
<ID>Q</ID>446 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>475</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>0.5,75</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>442 </input>
<input>
<ID>IN_2</ID>444 </input>
<input>
<ID>IN_3</ID>443 </input>
<input>
<ID>IN_4</ID>445 </input>
<input>
<ID>IN_5</ID>446 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>476</ID>
<type>AA_AND2</type>
<position>-198,173</position>
<input>
<ID>IN_0</ID>424 </input>
<input>
<ID>IN_1</ID>426 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>477</ID>
<type>AA_AND2</type>
<position>370,-1520</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>AA_AND2</type>
<position>-69.5,100</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>479</ID>
<type>AA_AND2</type>
<position>-52.5,99</position>
<input>
<ID>IN_0</ID>437 </input>
<input>
<ID>IN_1</ID>444 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_AND2</type>
<position>-181,172</position>
<input>
<ID>IN_0</ID>420 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>421 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>481</ID>
<type>AA_AND2</type>
<position>-37.5,98</position>
<input>
<ID>IN_0</ID>438 </input>
<input>
<ID>IN_1</ID>443 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>482</ID>
<type>AA_AND2</type>
<position>-20,97</position>
<input>
<ID>IN_0</ID>439 </input>
<input>
<ID>IN_1</ID>445 </input>
<output>
<ID>OUT</ID>440 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>483</ID>
<type>AA_AND2</type>
<position>-166,171</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>484</ID>
<type>BA_NAND4</type>
<position>2,100</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>443 </input>
<input>
<ID>IN_2</ID>445 </input>
<input>
<ID>IN_3</ID>446 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>485</ID>
<type>AE_DFF_LOW</type>
<position>-81,54.5</position>
<input>
<ID>IN_0</ID>441 </input>
<output>
<ID>OUT_0</ID>447 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>486</ID>
<type>AA_AND2</type>
<position>-148.5,170</position>
<input>
<ID>IN_0</ID>422 </input>
<input>
<ID>IN_1</ID>429 </input>
<output>
<ID>OUT</ID>423 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_DFF_LOW</type>
<position>-64.5,54.5</position>
<input>
<ID>IN_0</ID>442 </input>
<output>
<ID>OUT_0</ID>448 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>488</ID>
<type>AE_DFF_LOW</type>
<position>-50,54.5</position>
<input>
<ID>IN_0</ID>444 </input>
<output>
<ID>OUT_0</ID>449 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>489</ID>
<type>BA_NAND4</type>
<position>-126.5,173</position>
<input>
<ID>IN_0</ID>428 </input>
<input>
<ID>IN_1</ID>427 </input>
<input>
<ID>IN_2</ID>429 </input>
<input>
<ID>IN_3</ID>430 </input>
<output>
<ID>OUT</ID>406 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>490</ID>
<type>AE_DFF_LOW</type>
<position>-33,54.5</position>
<input>
<ID>IN_0</ID>443 </input>
<output>
<ID>OUT_0</ID>450 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>491</ID>
<type>AE_DFF_LOW</type>
<position>-17,54.5</position>
<input>
<ID>IN_0</ID>445 </input>
<output>
<ID>OUT_0</ID>451 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>492</ID>
<type>AE_DFF_LOW</type>
<position>1,54.5</position>
<input>
<ID>IN_0</ID>446 </input>
<output>
<ID>OUT_0</ID>452 </output>
<input>
<ID>clear</ID>401 </input>
<input>
<ID>clock</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>493</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>21,45</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>448 </input>
<input>
<ID>IN_2</ID>449 </input>
<input>
<ID>IN_3</ID>450 </input>
<input>
<ID>IN_4</ID>451 </input>
<input>
<ID>IN_5</ID>452 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_INVERTER</type>
<position>-91.5,147.5</position>
<input>
<ID>IN_0</ID>405 </input>
<output>
<ID>OUT_0</ID>454 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>495</ID>
<type>AE_DFF_LOW</type>
<position>-209.5,127.5</position>
<input>
<ID>IN_0</ID>424 </input>
<output>
<ID>OUT_0</ID>431 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>499</ID>
<type>AE_DFF_LOW</type>
<position>-193,127.5</position>
<input>
<ID>IN_0</ID>426 </input>
<output>
<ID>OUT_0</ID>432 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>500</ID>
<type>AE_DFF_LOW</type>
<position>-178.5,127.5</position>
<input>
<ID>IN_0</ID>428 </input>
<output>
<ID>OUT_0</ID>433 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>503</ID>
<type>AE_DFF_LOW</type>
<position>-161.5,127.5</position>
<input>
<ID>IN_0</ID>427 </input>
<output>
<ID>OUT_0</ID>434 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>505</ID>
<type>AE_DFF_LOW</type>
<position>-145.5,127.5</position>
<input>
<ID>IN_0</ID>429 </input>
<output>
<ID>OUT_0</ID>435 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>507</ID>
<type>AE_DFF_LOW</type>
<position>-127.5,127.5</position>
<input>
<ID>IN_0</ID>430 </input>
<output>
<ID>OUT_0</ID>436 </output>
<input>
<ID>clear</ID>405 </input>
<input>
<ID>clock</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>509</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-107.5,118</position>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_2</ID>433 </input>
<input>
<ID>IN_3</ID>434 </input>
<input>
<ID>IN_4</ID>435 </input>
<input>
<ID>IN_5</ID>436 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_AND2</type>
<position>-245,158.5</position>
<input>
<ID>IN_0</ID>1576 </input>
<input>
<ID>IN_1</ID>335 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>AE_DFF_LOW</type>
<position>-301,-8.5</position>
<input>
<ID>IN_0</ID>330 </input>
<output>
<ID>OUTINV_0</ID>336 </output>
<output>
<ID>OUT_0</ID>334 </output>
<input>
<ID>clock</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_TOGGLE</type>
<position>-313.5,-6.5</position>
<output>
<ID>OUT_0</ID>330 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>513</ID>
<type>AI_XOR2</type>
<position>243.5,-228.5</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>471 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AI_XOR2</type>
<position>257,-228.5</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>308 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_AND2</type>
<position>-284.5,2.5</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>333 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AI_XOR2</type>
<position>270,-228.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>475 </input>
<output>
<ID>OUT</ID>309 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>517</ID>
<type>AA_LABEL</type>
<position>-317.5,3</position>
<gparam>LABEL_TEXT On/Off Switch</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>518</ID>
<type>AI_XOR2</type>
<position>283,-228.5</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>477 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>519</ID>
<type>AI_XOR2</type>
<position>295.5,-229</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>311 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>AE_SMALL_INVERTER</type>
<position>-290.5,-9.5</position>
<input>
<ID>IN_0</ID>336 </input>
<output>
<ID>OUT_0</ID>337 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>521</ID>
<type>AI_XOR2</type>
<position>308,-229</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>481 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_LABEL</type>
<position>-162.5,-19</position>
<gparam>LABEL_TEXT Default Power</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>523</ID>
<type>AE_DFF_LOW</type>
<position>-251,-10.5</position>
<input>
<ID>IN_0</ID>331 </input>
<output>
<ID>OUTINV_0</ID>333 </output>
<output>
<ID>OUT_0</ID>389 </output>
<input>
<ID>clear</ID>337 </input>
<input>
<ID>clock</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>524</ID>
<type>BB_CLOCK</type>
<position>-266,-14</position>
<output>
<ID>CLK</ID>332 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>525</ID>
<type>AA_AND2</type>
<position>330.5,-1150.5</position>
<input>
<ID>IN_0</ID>459 </input>
<input>
<ID>IN_1</ID>458 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>526</ID>
<type>AA_TOGGLE</type>
<position>123.5,-279.5</position>
<output>
<ID>OUT_0</ID>2141 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND2</type>
<position>308,-1173.5</position>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>460 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>AA_AND2</type>
<position>154.5,-346</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>482 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>529</ID>
<type>AA_AND2</type>
<position>154,-337.5</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>530</ID>
<type>AA_AND2</type>
<position>153.5,-329</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>AA_AND2</type>
<position>153,-321</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>532</ID>
<type>AA_AND2</type>
<position>152.5,-312.5</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>533</ID>
<type>AA_AND2</type>
<position>152.5,-304</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>603 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>534</ID>
<type>AI_XOR2</type>
<position>265,-1118.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>465 </input>
<output>
<ID>OUT</ID>297 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>535</ID>
<type>AA_LABEL</type>
<position>116.5,-119.5</position>
<gparam>LABEL_TEXT Zone 1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>536</ID>
<type>AI_XOR2</type>
<position>278.5,-1118.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>298 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_LABEL</type>
<position>124,-269</position>
<gparam>LABEL_TEXT Zone 2</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>538</ID>
<type>AI_XOR2</type>
<position>291.5,-1118.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>469 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>539</ID>
<type>AI_XOR2</type>
<position>304.5,-1118.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>484 </input>
<output>
<ID>OUT</ID>302 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>540</ID>
<type>AI_XOR2</type>
<position>317,-1119</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>486 </input>
<output>
<ID>OUT</ID>303 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>542</ID>
<type>AI_XOR2</type>
<position>329.5,-1119</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>488 </input>
<output>
<ID>OUT</ID>305 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>543</ID>
<type>BE_JKFF_LOW_NT</type>
<position>222.5,-191.5</position>
<input>
<ID>J</ID>470 </input>
<output>
<ID>Q</ID>471 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>544</ID>
<type>AI_XOR2</type>
<position>356,-1629</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>545</ID>
<type>AA_LABEL</type>
<position>132,-989</position>
<gparam>LABEL_TEXT Zone 6</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>546</ID>
<type>BE_JKFF_LOW_NT</type>
<position>209.5,-181.5</position>
<input>
<ID>J</ID>472 </input>
<output>
<ID>Q</ID>473 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>547</ID>
<type>BE_JKFF_LOW_NT</type>
<position>196.5,-170.5</position>
<input>
<ID>J</ID>474 </input>
<output>
<ID>Q</ID>475 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>548</ID>
<type>BE_JKFF_LOW_NT</type>
<position>189,-161.5</position>
<input>
<ID>J</ID>476 </input>
<output>
<ID>Q</ID>477 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>549</ID>
<type>BE_JKFF_LOW_NT</type>
<position>180.5,-154</position>
<input>
<ID>J</ID>478 </input>
<output>
<ID>Q</ID>479 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>550</ID>
<type>BE_JKFF_LOW_NT</type>
<position>171.5,-146.5</position>
<input>
<ID>J</ID>480 </input>
<output>
<ID>Q</ID>481 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>551</ID>
<type>BE_JKFF_LOW_NT</type>
<position>212.5,-348</position>
<input>
<ID>J</ID>482 </input>
<output>
<ID>Q</ID>594 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2090</ID>
<type>BE_JKFF_LOW_NT</type>
<position>314.5,-293</position>
<input>
<ID>J</ID>1411 </input>
<output>
<ID>Q</ID>27 </output>
<input>
<ID>clear</ID>1577 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>552</ID>
<type>BE_JKFF_LOW_NT</type>
<position>204.5,-339.5</position>
<input>
<ID>J</ID>595 </input>
<output>
<ID>Q</ID>596 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>553</ID>
<type>BE_JKFF_LOW_NT</type>
<position>197.5,-331</position>
<input>
<ID>J</ID>597 </input>
<output>
<ID>Q</ID>598 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>554</ID>
<type>BE_JKFF_LOW_NT</type>
<position>188.5,-323</position>
<input>
<ID>J</ID>599 </input>
<output>
<ID>Q</ID>600 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2092</ID>
<type>AA_AND2</type>
<position>332.5,-297.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>461 </input>
<output>
<ID>OUT</ID>1835 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>BE_JKFF_LOW_NT</type>
<position>181.5,-314.5</position>
<input>
<ID>J</ID>601 </input>
<output>
<ID>Q</ID>602 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>556</ID>
<type>BE_JKFF_LOW_NT</type>
<position>173.5,-306</position>
<input>
<ID>J</ID>603 </input>
<output>
<ID>Q</ID>604 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2094</ID>
<type>AA_AND2</type>
<position>331.5,-348</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>1835 </input>
<output>
<ID>OUT</ID>1836 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>558</ID>
<type>BE_JKFF_LOW_NT</type>
<position>244,-1081.5</position>
<input>
<ID>J</ID>464 </input>
<output>
<ID>Q</ID>465 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2096</ID>
<type>AA_AND2</type>
<position>345,-345</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>1835 </input>
<output>
<ID>OUT</ID>1837 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>559</ID>
<type>BE_JKFF_LOW_NT</type>
<position>231,-1071.5</position>
<input>
<ID>J</ID>466 </input>
<output>
<ID>Q</ID>467 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>560</ID>
<type>BE_JKFF_LOW_NT</type>
<position>218,-1060.5</position>
<input>
<ID>J</ID>468 </input>
<output>
<ID>Q</ID>469 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2098</ID>
<type>AA_AND2</type>
<position>344.5,-337.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>1835 </input>
<output>
<ID>OUT</ID>1838 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>561</ID>
<type>AI_XOR2</type>
<position>321.5,-1166.5</position>
<input>
<ID>IN_0</ID>460 </input>
<input>
<ID>IN_1</ID>462 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2100</ID>
<type>AA_AND2</type>
<position>345.5,-329.5</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>1835 </input>
<output>
<ID>OUT</ID>1839 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>563</ID>
<type>BE_JKFF_LOW_NT</type>
<position>210.5,-1051.5</position>
<input>
<ID>J</ID>483 </input>
<output>
<ID>Q</ID>484 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2102</ID>
<type>AA_AND2</type>
<position>345.5,-323.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>1835 </input>
<output>
<ID>OUT</ID>1840 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>565</ID>
<type>BE_JKFF_LOW_NT</type>
<position>202,-1044</position>
<input>
<ID>J</ID>485 </input>
<output>
<ID>Q</ID>486 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>566</ID>
<type>CC_PULSE</type>
<position>165.5,-294</position>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2104</ID>
<type>AA_AND2</type>
<position>346,-318</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>1835 </input>
<output>
<ID>OUT</ID>1841 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>567</ID>
<type>BE_JKFF_LOW_NT</type>
<position>193,-1036.5</position>
<input>
<ID>J</ID>487 </input>
<output>
<ID>Q</ID>488 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2106</ID>
<type>AI_XOR2</type>
<position>353.5,-401.5</position>
<input>
<ID>IN_0</ID>1842 </input>
<input>
<ID>IN_1</ID>1843 </input>
<output>
<ID>OUT</ID>1844 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>568</ID>
<type>CC_PULSE</type>
<position>163,-138.5</position>
<output>
<ID>OUT_0</ID>609 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>569</ID>
<type>CC_PULSE</type>
<position>185,-1028.5</position>
<output>
<ID>OUT_0</ID>489 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>2108</ID>
<type>BA_NAND2</type>
<position>468,-268.5</position>
<input>
<ID>IN_0</ID>1844 </input>
<input>
<ID>IN_1</ID>1843 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>571</ID>
<type>AA_AND2</type>
<position>179,-1079.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>464 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_TOGGLE</type>
<position>326,-114.5</position>
<output>
<ID>OUT_0</ID>611 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>573</ID>
<type>AA_AND2</type>
<position>178.5,-1069.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>574</ID>
<type>AA_AND2</type>
<position>177,-1058.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>575</ID>
<type>AA_AND2</type>
<position>176.5,-1049.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>576</ID>
<type>AA_AND2</type>
<position>175.5,-1042</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>577</ID>
<type>AA_AND2</type>
<position>174.5,-1034.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>AE_DFF_LOW</type>
<position>269,-1127</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>306 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>579</ID>
<type>AE_DFF_LOW</type>
<position>287,-1361.5</position>
<input>
<ID>IN_0</ID>494 </input>
<output>
<ID>OUT_0</ID>500 </output>
<input>
<ID>clear</ID>165 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>580</ID>
<type>AE_DFF_LOW</type>
<position>300.5,-1361.5</position>
<input>
<ID>IN_0</ID>495 </input>
<output>
<ID>OUT_0</ID>501 </output>
<input>
<ID>clear</ID>165 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>581</ID>
<type>AE_DFF_LOW</type>
<position>315.5,-1361.5</position>
<input>
<ID>IN_0</ID>496 </input>
<output>
<ID>OUT_0</ID>502 </output>
<input>
<ID>clear</ID>165 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>582</ID>
<type>AE_DFF_LOW</type>
<position>326,-1361.5</position>
<input>
<ID>IN_0</ID>497 </input>
<output>
<ID>OUT_0</ID>503 </output>
<input>
<ID>clear</ID>165 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>583</ID>
<type>AE_DFF_LOW</type>
<position>339,-1361.5</position>
<input>
<ID>IN_0</ID>498 </input>
<output>
<ID>OUT_0</ID>504 </output>
<input>
<ID>clear</ID>165 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>584</ID>
<type>AE_SMALL_INVERTER</type>
<position>278,-1369</position>
<input>
<ID>IN_0</ID>499 </input>
<output>
<ID>OUT_0</ID>505 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>585</ID>
<type>AE_SMALL_INVERTER</type>
<position>293,-1369</position>
<input>
<ID>IN_0</ID>500 </input>
<output>
<ID>OUT_0</ID>506 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>586</ID>
<type>AE_SMALL_INVERTER</type>
<position>308,-1369</position>
<input>
<ID>IN_0</ID>501 </input>
<output>
<ID>OUT_0</ID>507 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>587</ID>
<type>AE_SMALL_INVERTER</type>
<position>319.5,-1368.5</position>
<input>
<ID>IN_0</ID>502 </input>
<output>
<ID>OUT_0</ID>508 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>588</ID>
<type>AE_SMALL_INVERTER</type>
<position>332.5,-1369</position>
<input>
<ID>IN_0</ID>503 </input>
<output>
<ID>OUT_0</ID>509 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>589</ID>
<type>AE_SMALL_INVERTER</type>
<position>345.5,-1368.5</position>
<input>
<ID>IN_0</ID>504 </input>
<output>
<ID>OUT_0</ID>510 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>591</ID>
<type>AA_AND4</type>
<position>296,-1385.5</position>
<input>
<ID>IN_0</ID>508 </input>
<input>
<ID>IN_1</ID>507 </input>
<input>
<ID>IN_2</ID>506 </input>
<input>
<ID>IN_3</ID>505 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>592</ID>
<type>AA_LABEL</type>
<position>186.5,-1255</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>593</ID>
<type>AA_AND2</type>
<position>332.5,-1384.5</position>
<input>
<ID>IN_0</ID>510 </input>
<input>
<ID>IN_1</ID>509 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>594</ID>
<type>AA_AND2</type>
<position>310,-1407.5</position>
<input>
<ID>IN_0</ID>512 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>595</ID>
<type>AI_XOR2</type>
<position>267,-1352.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>596</ID>
<type>AI_XOR2</type>
<position>280.5,-1352.5</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>517 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>597</ID>
<type>AI_XOR2</type>
<position>293.5,-1352.5</position>
<input>
<ID>IN_0</ID>1570 </input>
<input>
<ID>IN_1</ID>519 </input>
<output>
<ID>OUT</ID>495 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>AI_XOR2</type>
<position>306.5,-1352.5</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>521 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>599</ID>
<type>AI_XOR2</type>
<position>319,-1353</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>523 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>600</ID>
<type>BA_NAND2</type>
<position>558,-270</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AI_XOR2</type>
<position>331.5,-1353</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>525 </input>
<output>
<ID>OUT</ID>498 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_LABEL</type>
<position>133.5,-1231</position>
<gparam>LABEL_TEXT Zone 7</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>604</ID>
<type>AA_AND4</type>
<position>538,-251</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<input>
<ID>IN_2</ID>237 </input>
<input>
<ID>IN_3</ID>238 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>605</ID>
<type>BE_JKFF_LOW_NT</type>
<position>246,-1315.5</position>
<input>
<ID>J</ID>514 </input>
<output>
<ID>Q</ID>515 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>606</ID>
<type>BE_JKFF_LOW_NT</type>
<position>233,-1305.5</position>
<input>
<ID>J</ID>516 </input>
<output>
<ID>Q</ID>517 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>607</ID>
<type>BE_JKFF_LOW_NT</type>
<position>220,-1294.5</position>
<input>
<ID>J</ID>518 </input>
<output>
<ID>Q</ID>519 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>608</ID>
<type>AI_XOR2</type>
<position>323.5,-1400.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>609</ID>
<type>BE_JKFF_LOW_NT</type>
<position>212.5,-1285.5</position>
<input>
<ID>J</ID>520 </input>
<output>
<ID>Q</ID>521 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>610</ID>
<type>BE_JKFF_LOW_NT</type>
<position>204,-1278</position>
<input>
<ID>J</ID>522 </input>
<output>
<ID>Q</ID>523 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>611</ID>
<type>BE_JKFF_LOW_NT</type>
<position>195,-1270.5</position>
<input>
<ID>J</ID>524 </input>
<output>
<ID>Q</ID>525 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>612</ID>
<type>CC_PULSE</type>
<position>187,-1262.5</position>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>614</ID>
<type>AA_AND2</type>
<position>181,-1313.5</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>514 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AA_AND2</type>
<position>180.5,-1303.5</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_AND2</type>
<position>179,-1292.5</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>617</ID>
<type>AA_AND2</type>
<position>178.5,-1283.5</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>AA_AND2</type>
<position>177.5,-1276</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>619</ID>
<type>AA_AND2</type>
<position>176.5,-1268.5</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>620</ID>
<type>AE_DFF_LOW</type>
<position>271,-1361</position>
<input>
<ID>IN_0</ID>493 </input>
<output>
<ID>OUT_0</ID>499 </output>
<input>
<ID>clear</ID>165 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>621</ID>
<type>AE_DFF_LOW</type>
<position>296,-1588.5</position>
<input>
<ID>IN_0</ID>531 </input>
<output>
<ID>OUT_0</ID>537 </output>
<input>
<ID>clear</ID>1569 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>622</ID>
<type>AE_DFF_LOW</type>
<position>309.5,-1588.5</position>
<input>
<ID>IN_0</ID>532 </input>
<output>
<ID>OUT_0</ID>538 </output>
<input>
<ID>clear</ID>1569 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>623</ID>
<type>AE_DFF_LOW</type>
<position>324.5,-1588.5</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>539 </output>
<input>
<ID>clear</ID>1569 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>624</ID>
<type>AE_DFF_LOW</type>
<position>335,-1588.5</position>
<input>
<ID>IN_0</ID>534 </input>
<output>
<ID>OUT_0</ID>540 </output>
<input>
<ID>clear</ID>1569 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>625</ID>
<type>AE_DFF_LOW</type>
<position>348,-1588.5</position>
<input>
<ID>IN_0</ID>535 </input>
<output>
<ID>OUT_0</ID>541 </output>
<input>
<ID>clear</ID>1569 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>626</ID>
<type>AE_SMALL_INVERTER</type>
<position>287,-1596</position>
<input>
<ID>IN_0</ID>536 </input>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>627</ID>
<type>AE_SMALL_INVERTER</type>
<position>302,-1596</position>
<input>
<ID>IN_0</ID>537 </input>
<output>
<ID>OUT_0</ID>543 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>628</ID>
<type>AE_SMALL_INVERTER</type>
<position>317,-1596</position>
<input>
<ID>IN_0</ID>538 </input>
<output>
<ID>OUT_0</ID>544 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>629</ID>
<type>AE_SMALL_INVERTER</type>
<position>328.5,-1595.5</position>
<input>
<ID>IN_0</ID>539 </input>
<output>
<ID>OUT_0</ID>545 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>630</ID>
<type>AE_SMALL_INVERTER</type>
<position>341.5,-1596</position>
<input>
<ID>IN_0</ID>540 </input>
<output>
<ID>OUT_0</ID>546 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>631</ID>
<type>AE_SMALL_INVERTER</type>
<position>354.5,-1595.5</position>
<input>
<ID>IN_0</ID>541 </input>
<output>
<ID>OUT_0</ID>547 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>633</ID>
<type>AA_AND4</type>
<position>305,-1612.5</position>
<input>
<ID>IN_0</ID>545 </input>
<input>
<ID>IN_1</ID>544 </input>
<input>
<ID>IN_2</ID>543 </input>
<input>
<ID>IN_3</ID>542 </input>
<output>
<ID>OUT</ID>548 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>634</ID>
<type>AA_LABEL</type>
<position>195.5,-1482</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>635</ID>
<type>AA_AND2</type>
<position>341.5,-1611.5</position>
<input>
<ID>IN_0</ID>547 </input>
<input>
<ID>IN_1</ID>546 </input>
<output>
<ID>OUT</ID>549 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>636</ID>
<type>AA_AND2</type>
<position>319,-1634.5</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>548 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>637</ID>
<type>AI_XOR2</type>
<position>276,-1579.5</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>552 </input>
<output>
<ID>OUT</ID>530 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>638</ID>
<type>AI_XOR2</type>
<position>289.5,-1579.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>554 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>639</ID>
<type>AI_XOR2</type>
<position>302.5,-1579.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>556 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>640</ID>
<type>AI_XOR2</type>
<position>315.5,-1579.5</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>558 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>AI_XOR2</type>
<position>328,-1580</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>560 </input>
<output>
<ID>OUT</ID>534 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>643</ID>
<type>AI_XOR2</type>
<position>340.5,-1580</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>562 </input>
<output>
<ID>OUT</ID>535 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>644</ID>
<type>AA_AND2</type>
<position>500,-229</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>645</ID>
<type>AA_LABEL</type>
<position>138.5,-1445</position>
<gparam>LABEL_TEXT Zone 8</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>647</ID>
<type>BE_JKFF_LOW_NT</type>
<position>255,-1542.5</position>
<input>
<ID>J</ID>551 </input>
<output>
<ID>Q</ID>552 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>648</ID>
<type>BE_JKFF_LOW_NT</type>
<position>242,-1532.5</position>
<input>
<ID>J</ID>553 </input>
<output>
<ID>Q</ID>554 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>649</ID>
<type>BE_JKFF_LOW_NT</type>
<position>229,-1521.5</position>
<input>
<ID>J</ID>555 </input>
<output>
<ID>Q</ID>556 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>650</ID>
<type>AI_XOR2</type>
<position>332.5,-1627.5</position>
<input>
<ID>IN_0</ID>548 </input>
<input>
<ID>IN_1</ID>549 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>651</ID>
<type>BE_JKFF_LOW_NT</type>
<position>221.5,-1512.5</position>
<input>
<ID>J</ID>557 </input>
<output>
<ID>Q</ID>558 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>652</ID>
<type>BE_JKFF_LOW_NT</type>
<position>213,-1505</position>
<input>
<ID>J</ID>559 </input>
<output>
<ID>Q</ID>560 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>653</ID>
<type>BE_JKFF_LOW_NT</type>
<position>204,-1497.5</position>
<input>
<ID>J</ID>561 </input>
<output>
<ID>Q</ID>562 </output>
<input>
<ID>clear</ID>611 </input>
<input>
<ID>clock</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>654</ID>
<type>CC_PULSE</type>
<position>196,-1489.5</position>
<output>
<ID>OUT_0</ID>563 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>656</ID>
<type>AA_AND2</type>
<position>190,-1540.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>551 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_AND2</type>
<position>189.5,-1530.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>658</ID>
<type>AA_AND2</type>
<position>188,-1519.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_AND2</type>
<position>187.5,-1510.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>557 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>660</ID>
<type>AA_AND2</type>
<position>186.5,-1503</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>559 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>661</ID>
<type>AA_AND2</type>
<position>185.5,-1495.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>561 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>662</ID>
<type>AE_DFF_LOW</type>
<position>280,-1588</position>
<input>
<ID>IN_0</ID>530 </input>
<output>
<ID>OUT_0</ID>536 </output>
<input>
<ID>clear</ID>1569 </input>
<input>
<ID>clock</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>664</ID>
<type>AA_LABEL</type>
<position>318.5,-107.5</position>
<gparam>LABEL_TEXT Reset Storage before saving</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>665</ID>
<type>AA_LABEL</type>
<position>240,-421</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-282,311.5,-270</points>
<intersection>-282 1</intersection>
<intersection>-270 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-282,320,-282</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,-270,311.5,-270</points>
<intersection>303 15</intersection>
<intersection>311.5 0</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>303,-276.5,303,-270</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<intersection>-270 2</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-414,315,-408</points>
<intersection>-414 2</intersection>
<intersection>-408 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308,-408,315,-408</points>
<connection>
<GID>7</GID>
<name>Q</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>315,-414,322,-414</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-566,316.5,-563.5</points>
<intersection>-566 2</intersection>
<intersection>-563.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-563.5,316.5,-563.5</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>316.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>316.5,-566,321,-566</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,-265.5,454,-260.5</points>
<connection>
<GID>1613</GID>
<name>OUT</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>470,-260.5,470,-255.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>454,-260.5,470,-260.5</points>
<intersection>454 0</intersection>
<intersection>470 1</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-399,335,-393.5</points>
<intersection>-399 2</intersection>
<intersection>-393.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331,-393.5,335,-393.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>335 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>335,-399,339,-399</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>335 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-496,337,-415</points>
<intersection>-496 2</intersection>
<intersection>-441.5 3</intersection>
<intersection>-415 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>328,-415,337,-415</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>337 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>336,-496,337,-496</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>337 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>337,-441.5,357.5,-441.5</points>
<intersection>337 0</intersection>
<intersection>357.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>357.5,-490.5,357.5,-441.5</points>
<intersection>-490.5 5</intersection>
<intersection>-482.5 6</intersection>
<intersection>-474.5 7</intersection>
<intersection>-464 8</intersection>
<intersection>-453 9</intersection>
<intersection>-441.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>351.5,-490.5,357.5,-490.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>357.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>352,-482.5,357.5,-482.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>357.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>353,-474.5,357.5,-474.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>357.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>353.5,-464,357.5,-464</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>357.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>353,-453,357.5,-453</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>357.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>320.5,-745.5,327.5,-745.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468,-265.5,468,-260.5</points>
<connection>
<GID>2108</GID>
<name>OUT</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>472,-260.5,472,-255.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>468,-260.5,472,-260.5</points>
<intersection>468 0</intersection>
<intersection>472 1</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>331,-944.5,335.5,-944.5</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-727.5,176,-725.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-727.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-727.5,180.5,-727.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>324.5,-1166.5,331,-1166.5</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>176,-721.5,194,-721.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>clear</name></connection>
<intersection>176 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>176,-721.5,176,-715.5</points>
<intersection>-721.5 1</intersection>
<intersection>-715.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>176,-715.5,191,-715.5</points>
<connection>
<GID>15</GID>
<name>J</name></connection>
<intersection>176 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>326.5,-1400.5,332.5,-1400.5</points>
<connection>
<GID>608</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197,-719.5,200,-719.5</points>
<connection>
<GID>15</GID>
<name>nQ</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>335.5,-1627.5,341.5,-1627.5</points>
<connection>
<GID>650</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254,-512.5,254,-497</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-497 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>254,-497,330,-497</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>254 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-512.5,267.5,-491.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-491.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-491.5,345.5,-491.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>267.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-512.5,280.5,-483.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-483.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280.5,-483.5,346,-483.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-568,133,-414.5</points>
<intersection>-568 13</intersection>
<intersection>-475.5 1</intersection>
<intersection>-465.5 3</intersection>
<intersection>-454.5 5</intersection>
<intersection>-445.5 7</intersection>
<intersection>-438 9</intersection>
<intersection>-430.5 11</intersection>
<intersection>-416 15</intersection>
<intersection>-414.5 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-475.5,164,-475.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133,-465.5,163.5,-465.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>133,-454.5,162,-454.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>133,-445.5,161.5,-445.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>133,-438,160.5,-438</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>133,-430.5,159.5,-430.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>133,-568,321,-568</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>133,-416,322,-416</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>119.5,-414.5,133,-414.5</points>
<connection>
<GID>1825</GID>
<name>OUT</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-512.5,293.5,-475.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-475.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293.5,-475.5,347,-475.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306,-513,306,-465</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-465 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306,-465,347.5,-465</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>306 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323.5,-296.5,323.5,-291</points>
<intersection>-296.5 2</intersection>
<intersection>-291 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-291,323.5,-291</points>
<connection>
<GID>2090</GID>
<name>Q</name></connection>
<intersection>323.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>323.5,-296.5,329.5,-296.5</points>
<connection>
<GID>2092</GID>
<name>IN_0</name></connection>
<intersection>323.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-513,318.5,-454</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-454 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-454,347,-454</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488.5,-573.5,488.5,-271.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>-573.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>296,-573.5,488.5,-573.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>296 5</intersection>
<intersection>334 4</intersection>
<intersection>488.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>334,-573.5,334,-569</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-573.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>296,-577,296,-573.5</points>
<intersection>-577 6</intersection>
<intersection>-573.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>296,-577,308,-577</points>
<connection>
<GID>55</GID>
<name>J</name></connection>
<intersection>296 5</intersection></hsegment></shape></wire>
<wire>
<ID>1568</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>227.5,-1620,262,-1620</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>262 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>262,-1620,262,-1619</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>-1620 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>487.5,-265.5,487.5,-260.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>474,-260.5,474,-255.5</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>474,-260.5,487.5,-260.5</points>
<intersection>474 1</intersection>
<intersection>487.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-1609,280,-1592</points>
<connection>
<GID>662</GID>
<name>clear</name></connection>
<intersection>-1609 1</intersection>
<intersection>-1592.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,-1609,280,-1609</points>
<connection>
<GID>177</GID>
<name>Q</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,-1592.5,348,-1592.5</points>
<connection>
<GID>625</GID>
<name>clear</name></connection>
<connection>
<GID>624</GID>
<name>clear</name></connection>
<connection>
<GID>623</GID>
<name>clear</name></connection>
<connection>
<GID>622</GID>
<name>clear</name></connection>
<connection>
<GID>621</GID>
<name>clear</name></connection>
<intersection>280 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>504,-266,504,-260.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>476,-260.5,476,-255.5</points>
<connection>
<GID>9</GID>
<name>IN_3</name></connection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>476,-260.5,504,-260.5</points>
<intersection>476 1</intersection>
<intersection>504 0</intersection></hsegment></shape></wire>
<wire>
<ID>1570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-1349.5,294.5,-1324.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>-1324.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,-1324.5,347,-1324.5</points>
<connection>
<GID>251</GID>
<name>OUT</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186.5,-726.5,221,-726.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>221 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>221,-726.5,221,-725.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>-726.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>327,-567,334,-567</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-252.5,247.5,-241</points>
<connection>
<GID>368</GID>
<name>clear</name></connection>
<intersection>-252.5 7</intersection>
<intersection>-241.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-241.5,315.5,-241.5</points>
<connection>
<GID>422</GID>
<name>clear</name></connection>
<connection>
<GID>415</GID>
<name>clear</name></connection>
<connection>
<GID>410</GID>
<name>clear</name></connection>
<connection>
<GID>403</GID>
<name>clear</name></connection>
<connection>
<GID>394</GID>
<name>clear</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>225,-252.5,247.5,-252.5</points>
<connection>
<GID>1783</GID>
<name>Q</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-248.5,172,-248.5,173</points>
<intersection>172 1</intersection>
<intersection>173 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-248.5,172,-244,172</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>-248.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-253.5,173,-248.5,173</points>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection>
<intersection>-248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-271,156,-262.5</points>
<intersection>-271 1</intersection>
<intersection>-262.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-271,158.5,-271</points>
<connection>
<GID>1785</GID>
<name>OUT</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-262.5,204,-262.5</points>
<connection>
<GID>1789</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>1574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-258.5,222,-258.5</points>
<connection>
<GID>1783</GID>
<name>clear</name></connection>
<connection>
<GID>1789</GID>
<name>OUT_0</name></connection>
<intersection>204 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>204,-258.5,204,-252.5</points>
<intersection>-258.5 1</intersection>
<intersection>-252.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>204,-252.5,219,-252.5</points>
<connection>
<GID>1783</GID>
<name>J</name></connection>
<intersection>204 3</intersection></hsegment></shape></wire>
<wire>
<ID>1575</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,-256.5,228,-256.5</points>
<connection>
<GID>1783</GID>
<name>nQ</name></connection>
<connection>
<GID>1791</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>1576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-237.5,162,-237.5,173</points>
<intersection>162 1</intersection>
<intersection>173 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-248,162,-237.5,162</points>
<intersection>-248 3</intersection>
<intersection>-237.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-238,173,-237.5,173</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<intersection>-237.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-248,159.5,-248,162</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>162 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,-562,347,-561</points>
<intersection>-562 1</intersection>
<intersection>-561 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,-562,486.5,-562</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<intersection>347 0</intersection>
<intersection>486.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-561,347,-561</points>
<intersection>341.5 6</intersection>
<intersection>347 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>486.5,-562,486.5,-271.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-562 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>341.5,-568,341.5,-561</points>
<intersection>-568 7</intersection>
<intersection>-561 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>340,-568,341.5,-568</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>341.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-297,196,-113</points>
<connection>
<GID>1793</GID>
<name>OUT_0</name></connection>
<intersection>-297 2</intersection>
<intersection>-266 1</intersection>
<intersection>-265 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-266,196,-266</points>
<connection>
<GID>1795</GID>
<name>IN_1</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>196,-297,314.5,-297</points>
<connection>
<GID>2090</GID>
<name>clear</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>196,-265,665.5,-265</points>
<intersection>196 0</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>665.5,-1616.5,665.5,-265</points>
<intersection>-1616.5 5</intersection>
<intersection>-1424.5 6</intersection>
<intersection>-1190 11</intersection>
<intersection>-965 15</intersection>
<intersection>-768.5 18</intersection>
<intersection>-583 21</intersection>
<intersection>-414 24</intersection>
<intersection>-265 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>268,-1616.5,665.5,-1616.5</points>
<intersection>268 10</intersection>
<intersection>665.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>249,-1424.5,665.5,-1424.5</points>
<connection>
<GID>267</GID>
<name>clear</name></connection>
<intersection>249 7</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>249,-1424.5,249,-1389.5</points>
<intersection>-1424.5 6</intersection>
<intersection>-1389.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>245.5,-1389.5,249,-1389.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>249 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>268,-1618,268,-1616.5</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>-1616.5 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>247,-1190,665.5,-1190</points>
<connection>
<GID>242</GID>
<name>clear</name></connection>
<intersection>247 12</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>247,-1190,247,-1156</points>
<intersection>-1190 11</intersection>
<intersection>-1156 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>243.5,-1156,247,-1156</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>247 12</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>248,-965,665.5,-965</points>
<connection>
<GID>188</GID>
<name>clear</name></connection>
<intersection>248 16</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>248,-965,248,-933</points>
<intersection>-965 15</intersection>
<intersection>-933 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>245,-933,248,-933</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>248 16</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>230.5,-768.5,665.5,-768.5</points>
<connection>
<GID>162</GID>
<name>clear</name></connection>
<intersection>230.5 19</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>230.5,-768.5,230.5,-724.5</points>
<intersection>-768.5 18</intersection>
<intersection>-724.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>227,-724.5,230.5,-724.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>230.5 19</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>231.5,-583,665.5,-583</points>
<connection>
<GID>55</GID>
<name>clear</name></connection>
<intersection>231.5 22</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>231.5,-583,231.5,-557</points>
<intersection>-583 21</intersection>
<intersection>-557 23</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>228,-557,231.5,-557</points>
<connection>
<GID>1813</GID>
<name>IN_1</name></connection>
<intersection>231.5 22</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>211,-414,665.5,-414</points>
<connection>
<GID>7</GID>
<name>clear</name></connection>
<intersection>211 25</intersection>
<intersection>665.5 4</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>211,-414,211,-388</points>
<intersection>-414 24</intersection>
<intersection>-388 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>164,-388,211,-388</points>
<connection>
<GID>1801</GID>
<name>IN_1</name></connection>
<intersection>211 25</intersection></hsegment></shape></wire>
<wire>
<ID>1578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>164.5,-270,167,-270</points>
<connection>
<GID>1785</GID>
<name>IN_1</name></connection>
<intersection>167 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>167,-270,167,-267</points>
<intersection>-270 1</intersection>
<intersection>-267 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>167,-267,169.5,-267</points>
<connection>
<GID>1795</GID>
<name>OUT</name></connection>
<intersection>167 3</intersection></hsegment></shape></wire>
<wire>
<ID>1579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-390,146,-390</points>
<connection>
<GID>1798</GID>
<name>IN_0</name></connection>
<connection>
<GID>1797</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-383,219,-383</points>
<connection>
<GID>1796</GID>
<name>clear</name></connection>
<intersection>142 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>142,-386,142,-377</points>
<connection>
<GID>1798</GID>
<name>OUT_0</name></connection>
<intersection>-383 1</intersection>
<intersection>-377 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>142,-377,216,-377</points>
<connection>
<GID>1796</GID>
<name>J</name></connection>
<intersection>142 3</intersection></hsegment></shape></wire>
<wire>
<ID>1581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-381,225,-381</points>
<connection>
<GID>1799</GID>
<name>N_in0</name></connection>
<connection>
<GID>1796</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-360,243,-356.5</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<intersection>-360 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-360,244,-360</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>1583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-389,158,-389</points>
<connection>
<GID>1797</GID>
<name>IN_1</name></connection>
<connection>
<GID>1801</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,-377,247,-366</points>
<connection>
<GID>334</GID>
<name>clear</name></connection>
<intersection>-377 1</intersection>
<intersection>-366.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-377,247,-377</points>
<connection>
<GID>1796</GID>
<name>Q</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>247,-366.5,315,-366.5</points>
<connection>
<GID>98</GID>
<name>clear</name></connection>
<connection>
<GID>97</GID>
<name>clear</name></connection>
<connection>
<GID>92</GID>
<name>clear</name></connection>
<connection>
<GID>88</GID>
<name>clear</name></connection>
<connection>
<GID>75</GID>
<name>clear</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-360.5,256.5,-356.5</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256.5,-360.5,260,-360.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>256.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-560,177,-558</points>
<connection>
<GID>1810</GID>
<name>IN_0</name></connection>
<intersection>-560 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-560,181.5,-560</points>
<connection>
<GID>1809</GID>
<name>OUT</name></connection>
<intersection>177 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-360.5,269.5,-356.5</points>
<connection>
<GID>330</GID>
<name>OUT</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,-360.5,273.5,-360.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1592</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-554,195,-554</points>
<connection>
<GID>1810</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1808</GID>
<name>clear</name></connection>
<intersection>177 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177,-554,177,-548</points>
<intersection>-554 1</intersection>
<intersection>-548 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177,-548,192,-548</points>
<connection>
<GID>1808</GID>
<name>J</name></connection>
<intersection>177 3</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-360.5,285.5,-356.5</points>
<intersection>-360.5 1</intersection>
<intersection>-356.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>285.5,-360.5,288.5,-360.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>282.5,-356.5,285.5,-356.5</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-552,201,-552</points>
<connection>
<GID>1808</GID>
<name>nQ</name></connection>
<connection>
<GID>1811</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-359,295,-357</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>-359 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295,-359,299,-359</points>
<intersection>295 0</intersection>
<intersection>299 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>299,-360.5,299,-359</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-359 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-359,307.5,-357</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<intersection>-359 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>307.5,-359,312,-359</points>
<intersection>307.5 0</intersection>
<intersection>312 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>312,-360.5,312,-359</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-359 1</intersection></vsegment></shape></wire>
<wire>
<ID>1595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>187.5,-559,222,-559</points>
<connection>
<GID>1809</GID>
<name>IN_1</name></connection>
<intersection>222 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>222,-559,222,-558</points>
<connection>
<GID>1813</GID>
<name>OUT</name></connection>
<intersection>-559 1</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254,-368,254,-360</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-360 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,-360,254,-360</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>254 0</intersection></hsegment></shape></wire>
<wire>
<ID>1596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-548,257,-528</points>
<connection>
<GID>147</GID>
<name>clear</name></connection>
<intersection>-548 1</intersection>
<intersection>-528.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-548,257,-548</points>
<connection>
<GID>1808</GID>
<name>Q</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257,-528.5,325,-528.5</points>
<connection>
<GID>33</GID>
<name>clear</name></connection>
<connection>
<GID>31</GID>
<name>clear</name></connection>
<connection>
<GID>27</GID>
<name>clear</name></connection>
<connection>
<GID>14</GID>
<name>clear</name></connection>
<connection>
<GID>1</GID>
<name>clear</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-368,269,-360.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-360.5,269,-360.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-368,284,-360.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,-360.5,284,-360.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-367.5,295.5,-360.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,-360.5,295.5,-360.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,-368,308.5,-360.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>305,-360.5,308.5,-360.5</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>308.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,-367.5,321.5,-360.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,-360.5,321.5,-360.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>321.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254,-377.5,254,-372</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>-377.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>269,-383.5,269,-377.5</points>
<connection>
<GID>325</GID>
<name>IN_3</name></connection>
<intersection>-377.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>254,-377.5,269,-377.5</points>
<intersection>254 0</intersection>
<intersection>269 1</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-377,269,-372</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-377 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>271,-383.5,271,-377</points>
<connection>
<GID>325</GID>
<name>IN_2</name></connection>
<intersection>-377 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>269,-377,271,-377</points>
<intersection>269 0</intersection>
<intersection>271 1</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-377.5,284,-372</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-377.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>273,-383.5,273,-377.5</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>-377.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>273,-377.5,284,-377.5</points>
<intersection>273 1</intersection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-378.5,295.5,-371.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>-378.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>275,-383.5,275,-378.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>-378.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>275,-378.5,295.5,-378.5</points>
<intersection>275 1</intersection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-582,320.5,-577</points>
<intersection>-582 2</intersection>
<intersection>-577 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-577,320.5,-577</points>
<connection>
<GID>55</GID>
<name>Q</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,-582,327.5,-582</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253,-522,253,-518.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>-522 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253,-522,254,-522</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>253 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-694.5,262,-679</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-679 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-679,332.5,-679</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,-678,339.5,-583</points>
<intersection>-678 2</intersection>
<intersection>-616 3</intersection>
<intersection>-583 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,-583,339.5,-583</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>338.5,-678,339.5,-678</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>339.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>339.5,-616,352.5,-616</points>
<intersection>339.5 0</intersection>
<intersection>352.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>352.5,-666,352.5,-616</points>
<intersection>-666 6</intersection>
<intersection>-657.5 5</intersection>
<intersection>-650 7</intersection>
<intersection>-641 8</intersection>
<intersection>-633 9</intersection>
<intersection>-616 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>348.5,-657.5,352.5,-657.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>352.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>348.5,-666,352.5,-666</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>352.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>349.5,-650,352.5,-650</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>352.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>350,-641,352.5,-641</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>352.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>350.5,-633,352.5,-633</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>352.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-522.5,266.5,-518.5</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-522.5,270,-522.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-522.5,279.5,-518.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,-522.5,283.5,-522.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-694.5,275.5,-667</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-667 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-667,342.5,-667</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>275.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,100,8.5,102.5</points>
<intersection>100 2</intersection>
<intersection>102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,102.5,12.5,102.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,100,8.5,100</points>
<connection>
<GID>484</GID>
<name>OUT</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-522.5,295.5,-518.5</points>
<intersection>-522.5 1</intersection>
<intersection>-518.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-522.5,298.5,-522.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>292.5,-518.5,295.5,-518.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305,-521,305,-519</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-521 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>305,-521,309,-521</points>
<intersection>305 0</intersection>
<intersection>309 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>309,-522.5,309,-521</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-521 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-521,317.5,-519</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-521 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-521,322,-521</points>
<intersection>317.5 0</intersection>
<intersection>322 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>322,-522.5,322,-521</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-521 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-530,264,-522</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-522 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-522,264,-522</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>264 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,-530,279,-522.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-522.5,279,-522.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>279 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-530,294,-522.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289.5,-522.5,294,-522.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,-529.5,305.5,-522.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,-522.5,305.5,-522.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>305.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-530,318.5,-522.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-522.5,318.5,-522.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,-529.5,331.5,-522.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-522.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>328,-522.5,331.5,-522.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>331.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-539.5,264,-534</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-539.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>279,-545.5,279,-539.5</points>
<connection>
<GID>74</GID>
<name>IN_3</name></connection>
<intersection>-539.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>264,-539.5,279,-539.5</points>
<intersection>264 0</intersection>
<intersection>279 1</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,-539,279,-534</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-539 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>281,-545.5,281,-539</points>
<connection>
<GID>74</GID>
<name>IN_2</name></connection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>279,-539,281,-539</points>
<intersection>279 0</intersection>
<intersection>281 1</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-694.5,288.5,-658.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-658.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-658.5,342.5,-658.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-539.5,294,-534</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-539.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>283,-545.5,283,-539.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-539.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>283,-539.5,294,-539.5</points>
<intersection>283 1</intersection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,-540.5,305.5,-533.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>-540.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>285,-545.5,285,-540.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-540.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>285,-540.5,305.5,-540.5</points>
<intersection>285 1</intersection>
<intersection>305.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-694.5,301.5,-651</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-651 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>301.5,-651,343.5,-651</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-539,318.5,-534</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-539 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>317.5,-544.5,317.5,-539</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>317.5,-539,318.5,-539</points>
<intersection>317.5 1</intersection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,-539,331.5,-533.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>-539 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>319.5,-544.5,319.5,-539</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-539 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>319.5,-539,331.5,-539</points>
<intersection>319.5 1</intersection>
<intersection>331.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-559,282,-551.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-559 9</intersection>
<intersection>-554.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>295,-567.5,295,-554.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>-562.5 7</intersection>
<intersection>-554.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>282,-554.5,295,-554.5</points>
<intersection>282 0</intersection>
<intersection>295 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>295,-562.5,306.5,-562.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>295 1</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>228,-559,282,-559</points>
<connection>
<GID>1813</GID>
<name>IN_0</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-554,318.5,-550.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>-554 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>297,-567.5,297,-554</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-564.5 6</intersection>
<intersection>-561 8</intersection>
<intersection>-554 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>297,-554,318.5,-554</points>
<intersection>297 1</intersection>
<intersection>318.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>297,-564.5,306.5,-564.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>297 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187.5,-561,297,-561</points>
<connection>
<GID>1809</GID>
<name>IN_0</name></connection>
<intersection>297 1</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-695,314,-642</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>-642 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-642,344,-642</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-695,326.5,-634</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-634 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326.5,-634,344.5,-634</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<intersection>326.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,-746.5,337.5,-746</points>
<intersection>-746.5 1</intersection>
<intersection>-746 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,-746.5,337.5,-746.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>337.5,-746,342,-746</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-476.5,229,-476.5</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252,-512.5,252,-476.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-476.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-476.5,252,-476.5</points>
<connection>
<GID>123</GID>
<name>Q</name></connection>
<intersection>252 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169.5,-466.5,216,-466.5</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<connection>
<GID>125</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-512.5,265.5,-466.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-466.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-466.5,265.5,-466.5</points>
<connection>
<GID>125</GID>
<name>Q</name></connection>
<intersection>265.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,-455.5,203,-455.5</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<connection>
<GID>126</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-512.5,278.5,-455.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>-455.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209,-455.5,278.5,-455.5</points>
<connection>
<GID>126</GID>
<name>Q</name></connection>
<intersection>278.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-446.5,195.5,-446.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-512.5,291.5,-446.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-446.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-446.5,291.5,-446.5</points>
<connection>
<GID>129</GID>
<name>Q</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166.5,-439,187,-439</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<connection>
<GID>130</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-513,304,-439</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>-439 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-439,304,-439</points>
<connection>
<GID>130</GID>
<name>Q</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165.5,-431.5,178,-431.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-513,316.5,-431.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-431.5,316.5,-431.5</points>
<connection>
<GID>134</GID>
<name>Q</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-478.5,173,-427.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>-478.5 7</intersection>
<intersection>-468.5 5</intersection>
<intersection>-457.5 8</intersection>
<intersection>-448.5 3</intersection>
<intersection>-441 9</intersection>
<intersection>-433.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,-433.5,178,-433.5</points>
<connection>
<GID>134</GID>
<name>clock</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>173,-448.5,195.5,-448.5</points>
<connection>
<GID>129</GID>
<name>clock</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>173,-468.5,216,-468.5</points>
<connection>
<GID>125</GID>
<name>clock</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>173,-478.5,229,-478.5</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>173,-457.5,203,-457.5</points>
<connection>
<GID>126</GID>
<name>clock</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>173,-441,187,-441</points>
<connection>
<GID>130</GID>
<name>clock</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-762.5,304,-755.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>-762.5 7</intersection>
<intersection>-756 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-756,505,-756</points>
<intersection>304 0</intersection>
<intersection>342 5</intersection>
<intersection>505 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>505,-756,505,-272</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>-756 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>342,-756,342,-748</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>-756 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>304,-762.5,316,-762.5</points>
<connection>
<GID>162</GID>
<name>J</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>348,-742,503,-742</points>
<intersection>348 11</intersection>
<intersection>364.5 12</intersection>
<intersection>503 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>503,-742,503,-272</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-742 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>348,-747,348,-742</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>-742 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>364.5,-747,364.5,-742</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<intersection>-742 1</intersection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265,-715.5,265,-710</points>
<connection>
<GID>278</GID>
<name>clear</name></connection>
<intersection>-715.5 1</intersection>
<intersection>-710.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,-715.5,265,-715.5</points>
<connection>
<GID>15</GID>
<name>Q</name></connection>
<intersection>265 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265,-710.5,333,-710.5</points>
<connection>
<GID>200</GID>
<name>clear</name></connection>
<connection>
<GID>199</GID>
<name>clear</name></connection>
<connection>
<GID>198</GID>
<name>clear</name></connection>
<connection>
<GID>197</GID>
<name>clear</name></connection>
<connection>
<GID>196</GID>
<name>clear</name></connection>
<intersection>265 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-936,194,-934</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-936 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,-936,198.5,-936</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>194 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,-930,212,-930</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>clear</name></connection>
<intersection>194 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>194,-930,194,-924</points>
<intersection>-930 1</intersection>
<intersection>-924 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>194,-924,209,-924</points>
<connection>
<GID>40</GID>
<name>J</name></connection>
<intersection>194 3</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-928,218,-928</points>
<connection>
<GID>47</GID>
<name>N_in0</name></connection>
<connection>
<GID>40</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204.5,-935,239,-935</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>239 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239,-935,239,-934</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>-935 1</intersection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-924,275.5,-909</points>
<connection>
<GID>320</GID>
<name>clear</name></connection>
<intersection>-924 1</intersection>
<intersection>-909.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215,-924,275.5,-924</points>
<connection>
<GID>40</GID>
<name>Q</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>275.5,-909.5,343.5,-909.5</points>
<connection>
<GID>283</GID>
<name>clear</name></connection>
<connection>
<GID>282</GID>
<name>clear</name></connection>
<connection>
<GID>281</GID>
<name>clear</name></connection>
<connection>
<GID>280</GID>
<name>clear</name></connection>
<connection>
<GID>279</GID>
<name>clear</name></connection>
<intersection>275.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-1159,192.5,-1157</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-1159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,-1159,197,-1159</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192.5,-1153,210.5,-1153</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>clear</name></connection>
<intersection>192.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>192.5,-1153,192.5,-1147</points>
<intersection>-1153 1</intersection>
<intersection>-1147 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>192.5,-1147,207.5,-1147</points>
<connection>
<GID>54</GID>
<name>J</name></connection>
<intersection>192.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>213.5,-1151,216.5,-1151</points>
<connection>
<GID>54</GID>
<name>nQ</name></connection>
<connection>
<GID>148</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,-1158,237.5,-1158</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>237.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>237.5,-1158,237.5,-1157</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>-1158 1</intersection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-1147,269,-1131</points>
<connection>
<GID>578</GID>
<name>clear</name></connection>
<intersection>-1147 1</intersection>
<intersection>-1131.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-1147,269,-1147</points>
<connection>
<GID>54</GID>
<name>Q</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269,-1131.5,337,-1131.5</points>
<connection>
<GID>335</GID>
<name>clear</name></connection>
<connection>
<GID>324</GID>
<name>clear</name></connection>
<connection>
<GID>323</GID>
<name>clear</name></connection>
<connection>
<GID>322</GID>
<name>clear</name></connection>
<connection>
<GID>321</GID>
<name>clear</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-1392.5,194.5,-1390.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-1392.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,-1392.5,199,-1392.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-1386.5,212.5,-1386.5</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<connection>
<GID>160</GID>
<name>clear</name></connection>
<intersection>194.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>194.5,-1386.5,194.5,-1380.5</points>
<intersection>-1386.5 1</intersection>
<intersection>-1380.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>194.5,-1380.5,209.5,-1380.5</points>
<connection>
<GID>160</GID>
<name>J</name></connection>
<intersection>194.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215.5,-1384.5,218.5,-1384.5</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-1391.5,239.5,-1391.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>239.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239.5,-1391.5,239.5,-1390.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>-1391.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-1380.5,271,-1365</points>
<connection>
<GID>620</GID>
<name>clear</name></connection>
<intersection>-1380.5 1</intersection>
<intersection>-1365.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-1380.5,271,-1380.5</points>
<connection>
<GID>160</GID>
<name>Q</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>271,-1365.5,339,-1365.5</points>
<connection>
<GID>583</GID>
<name>clear</name></connection>
<connection>
<GID>582</GID>
<name>clear</name></connection>
<connection>
<GID>581</GID>
<name>clear</name></connection>
<connection>
<GID>580</GID>
<name>clear</name></connection>
<connection>
<GID>579</GID>
<name>clear</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-1621,217,-1619</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-1621 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,-1621,221.5,-1621</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-1615,235,-1615</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<connection>
<GID>177</GID>
<name>clear</name></connection>
<intersection>217 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>217,-1615,217,-1609</points>
<intersection>-1615 1</intersection>
<intersection>-1609 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>217,-1609,232,-1609</points>
<connection>
<GID>177</GID>
<name>J</name></connection>
<intersection>217 3</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238,-1613,241,-1613</points>
<connection>
<GID>177</GID>
<name>nQ</name></connection>
<connection>
<GID>183</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323.5,-773,323.5,-762.5</points>
<intersection>-773 2</intersection>
<intersection>-762.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-762.5,323.5,-762.5</points>
<connection>
<GID>162</GID>
<name>Q</name></connection>
<intersection>323.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>323.5,-773,325.5,-773</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>323.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-893.5,272.5,-845.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>-845.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272.5,-845.5,345,-845.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>272.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>353,-844.5,353,-774</points>
<intersection>-844.5 2</intersection>
<intersection>-797.5 3</intersection>
<intersection>-774 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331.5,-774,353,-774</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-844.5,353,-844.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>353 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>353,-797.5,370.5,-797.5</points>
<intersection>353 0</intersection>
<intersection>365.5 9</intersection>
<intersection>370.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>370.5,-836,370.5,-797.5</points>
<intersection>-836 5</intersection>
<intersection>-826 6</intersection>
<intersection>-819 7</intersection>
<intersection>-809.5 8</intersection>
<intersection>-797.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>363,-836,370.5,-836</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>370.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>363,-826,370.5,-826</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>370.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>364.5,-819,370.5,-819</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>370.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>365,-809.5,370.5,-809.5</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>370.5 4</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>365.5,-802.5,365.5,-797.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>-797.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-893.5,286,-834</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>-834 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-834,357,-834</points>
<intersection>286 0</intersection>
<intersection>357 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>357,-837,357,-834</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>-834 1</intersection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299,-893.5,299,-825.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-825.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>299,-825.5,357,-825.5</points>
<intersection>299 0</intersection>
<intersection>357 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>357,-827,357,-825.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>-825.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-893.5,312,-818</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-818 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312,-818,358.5,-818</points>
<intersection>312 0</intersection>
<intersection>358.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>358.5,-820,358.5,-818</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<intersection>-818 1</intersection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,-894,324.5,-810.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-810.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324.5,-810.5,359,-810.5</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-894,337,-803.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-803.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>337,-803.5,359.5,-803.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>337 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,-945.5,344,-945</points>
<intersection>-945.5 1</intersection>
<intersection>-945 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>341.5,-945.5,344,-945.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>344 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>344,-945,347,-945</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>344 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314.5,-959,314.5,-954.5</points>
<connection>
<GID>294</GID>
<name>OUT</name></connection>
<intersection>-959 7</intersection>
<intersection>-955 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314.5,-955,520,-955</points>
<intersection>314.5 0</intersection>
<intersection>347 5</intersection>
<intersection>520 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>520,-955,520,-272.5</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>-955 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>347,-955,347,-947</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>-955 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>314.5,-959,324,-959</points>
<connection>
<GID>188</GID>
<name>J</name></connection>
<intersection>314.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>358,-946,358,-945.5</points>
<intersection>-946 2</intersection>
<intersection>-945.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358,-945.5,518,-945.5</points>
<connection>
<GID>184</GID>
<name>N_in0</name></connection>
<intersection>358 0</intersection>
<intersection>518 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353,-946,358,-946</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>358 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>518,-945.5,518,-272.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>-945.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>334,-968.5,334,-959</points>
<intersection>-968.5 2</intersection>
<intersection>-959 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330,-959,334,-959</points>
<connection>
<GID>188</GID>
<name>Q</name></connection>
<intersection>334 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>334,-968.5,338.5,-968.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>334 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343,-1103,343,-969.5</points>
<intersection>-1103 2</intersection>
<intersection>-1045.5 3</intersection>
<intersection>-969.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>343,-969.5,344.5,-969.5</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>343 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,-1103,343,-1103</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>343 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>343,-1045.5,362,-1045.5</points>
<intersection>343 0</intersection>
<intersection>362 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>362,-1097,362,-1045.5</points>
<intersection>-1097 5</intersection>
<intersection>-1087.5 6</intersection>
<intersection>-1078 7</intersection>
<intersection>-1069.5 8</intersection>
<intersection>-1061 9</intersection>
<intersection>-1045.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>353,-1097,362,-1097</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>362 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>353,-1087.5,362,-1087.5</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>362 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>354,-1078,362,-1078</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>362 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>354.5,-1069.5,362,-1069.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>362 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>355.5,-1061,362,-1061</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>362 4</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-1115.5,266,-1104</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>-1104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-1104,336,-1104</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>266 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-747.5,141,-584</points>
<intersection>-747.5 13</intersection>
<intersection>-657.5 1</intersection>
<intersection>-647.5 3</intersection>
<intersection>-636.5 5</intersection>
<intersection>-627.5 7</intersection>
<intersection>-620 9</intersection>
<intersection>-612.5 11</intersection>
<intersection>-591.5 16</intersection>
<intersection>-584 15</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-657.5,172,-657.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>141,-647.5,171.5,-647.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>141,-636.5,170,-636.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>141,-627.5,169.5,-627.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>141,-620,168.5,-620</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>141,-612.5,167.5,-612.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>141,-747.5,327.5,-747.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>141,-584,327.5,-584</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>133,-591.5,141,-591.5</points>
<intersection>133 17</intersection>
<intersection>141 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>133,-591.5,133,-591</points>
<connection>
<GID>1829</GID>
<name>OUT</name></connection>
<intersection>-591.5 16</intersection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-704,261,-700.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>-704 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261,-704,262,-704</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>261 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-704.5,274.5,-700.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274.5,-704.5,278,-704.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-704.5,287.5,-700.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-704.5,291.5,-704.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>287.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-704.5,303.5,-700.5</points>
<intersection>-704.5 1</intersection>
<intersection>-700.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-704.5,306.5,-704.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>303.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>300.5,-700.5,303.5,-700.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-703,313,-701</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<intersection>-703 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-703,317,-703</points>
<intersection>313 0</intersection>
<intersection>317 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>317,-704.5,317,-703</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-703 1</intersection></vsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,-703,325.5,-701</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>-703 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325.5,-703,330,-703</points>
<intersection>325.5 0</intersection>
<intersection>330 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>330,-704.5,330,-703</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>-703 1</intersection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-712,272,-704</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-704 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,-704,272,-704</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<intersection>272 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-712,287,-704.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284,-704.5,287,-704.5</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>287 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-712,302,-704.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297.5,-704.5,302,-704.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-711.5,313.5,-704.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-704.5,313.5,-704.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-712,326.5,-704.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,-704.5,326.5,-704.5</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>326.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,-711.5,339.5,-704.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-704.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,-704.5,339.5,-704.5</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-721.5,272,-716</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>-721.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>287,-727.5,287,-721.5</points>
<connection>
<GID>208</GID>
<name>IN_3</name></connection>
<intersection>-721.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>272,-721.5,287,-721.5</points>
<intersection>272 0</intersection>
<intersection>287 1</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-721,287,-716</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>-721 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>289,-727.5,289,-721</points>
<connection>
<GID>208</GID>
<name>IN_2</name></connection>
<intersection>-721 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>287,-721,289,-721</points>
<intersection>287 0</intersection>
<intersection>289 1</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-721.5,302,-716</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-721.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>291,-727.5,291,-721.5</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>-721.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291,-721.5,302,-721.5</points>
<intersection>291 1</intersection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-722.5,313.5,-715.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>-722.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>293,-727.5,293,-722.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-722.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>293,-722.5,313.5,-722.5</points>
<intersection>293 1</intersection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-721,326.5,-716</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<intersection>-721 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>325.5,-726.5,325.5,-721</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>-721 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>325.5,-721,326.5,-721</points>
<intersection>325.5 1</intersection>
<intersection>326.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,-721,339.5,-715.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>-721 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>327.5,-726.5,327.5,-721</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>-721 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>327.5,-721,339.5,-721</points>
<intersection>327.5 1</intersection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-736.5,290,-733.5</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>-736.5 2</intersection>
<intersection>-734 8</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>303,-749.5,303,-736.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>-744.5 7</intersection>
<intersection>-736.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290,-736.5,303,-736.5</points>
<intersection>290 0</intersection>
<intersection>303 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>303,-744.5,314.5,-744.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>303 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>227,-734,290,-734</points>
<intersection>227 9</intersection>
<intersection>290 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>227,-734,227,-726.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-734 8</intersection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-1115.5,279.5,-1098</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>-1098 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,-1098,347,-1098</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-1115.5,292.5,-1088.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>-1088.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-1088.5,347,-1088.5</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,-1115.5,305.5,-1079</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>-1079 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>305.5,-1079,348,-1079</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>305.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318,-1116,318,-1070.5</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>-1070.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,-1070.5,348.5,-1070.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>318 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-736,326.5,-732.5</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>-736 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>305,-749.5,305,-736</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-746.5 6</intersection>
<intersection>-740 7</intersection>
<intersection>-736 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>305,-736,326.5,-736</points>
<intersection>305 1</intersection>
<intersection>326.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>305,-746.5,314.5,-746.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>305 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>186.5,-740,305,-740</points>
<intersection>186.5 8</intersection>
<intersection>305 1</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>186.5,-740,186.5,-728.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-740 7</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,-1116,330.5,-1062</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>-1062 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>330.5,-1062,349.5,-1062</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<intersection>330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>337,-1167.5,343.5,-1167.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-1184,308,-1176.5</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<intersection>-1184 4</intersection>
<intersection>-1177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308,-1177.5,534,-1177.5</points>
<intersection>308 0</intersection>
<intersection>343.5 7</intersection>
<intersection>534 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>534,-1177.5,534,-272.5</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>-1177.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>308,-1184,318.5,-1184</points>
<connection>
<GID>242</GID>
<name>J</name></connection>
<intersection>308 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>343.5,-1177.5,343.5,-1169.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>-1177.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-1168.5,354.5,-1167.5</points>
<intersection>-1168.5 2</intersection>
<intersection>-1167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354.5,-1167.5,532,-1167.5</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>354.5 0</intersection>
<intersection>532 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-1168.5,354.5,-1168.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>354.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>532,-1167.5,532,-272.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>-1167.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-1186.5,328.5,-1184</points>
<intersection>-1186.5 2</intersection>
<intersection>-1184 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324.5,-1184,328.5,-1184</points>
<connection>
<GID>242</GID>
<name>Q</name></connection>
<intersection>328.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>328.5,-1186.5,332.5,-1186.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268,-1349.5,268,-1343.5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>-1343.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,-1343.5,336.5,-1343.5</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<intersection>268 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343.5,-1342.5,343.5,-1187.5</points>
<intersection>-1342.5 2</intersection>
<intersection>-1279.5 3</intersection>
<intersection>-1187.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338.5,-1187.5,343.5,-1187.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342.5,-1342.5,343.5,-1342.5</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<intersection>343.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>343.5,-1279.5,364,-1279.5</points>
<intersection>343.5 0</intersection>
<intersection>364 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>364,-1333,364,-1279.5</points>
<intersection>-1333 5</intersection>
<intersection>-1323.5 11</intersection>
<intersection>-1315 13</intersection>
<intersection>-1306.5 15</intersection>
<intersection>-1299 17</intersection>
<intersection>-1279.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>353.5,-1333,364,-1333</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>364 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>353,-1323.5,364,-1323.5</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>364 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>353.5,-1315,364,-1315</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>364 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>353.5,-1306.5,364,-1306.5</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>364 4</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>354,-1299,364,-1299</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>364 4</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-1349.5,281.5,-1334</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>-1334 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-1334,347.5,-1334</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-1349.5,307.5,-1316</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>-1316 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>307.5,-1316,347.5,-1316</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>307.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-1350,320,-1307.5</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>-1307.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-1307.5,347.5,-1307.5</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-1350,332.5,-1300</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>-1300 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332.5,-1300,348,-1300</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>332.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-1401.5,341.5,-1400.5</points>
<intersection>-1401.5 1</intersection>
<intersection>-1400.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338.5,-1401.5,341.5,-1401.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341.5,-1400.5,345,-1400.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-1418.5,310,-1410.5</points>
<connection>
<GID>594</GID>
<name>OUT</name></connection>
<intersection>-1418.5 8</intersection>
<intersection>-1412 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-1412,547,-1412</points>
<intersection>310 0</intersection>
<intersection>344.5 5</intersection>
<intersection>547 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>547,-1412,547,-272.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>-1412 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>344.5,-1412,344.5,-1402.5</points>
<intersection>-1412 1</intersection>
<intersection>-1402.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>344.5,-1402.5,345,-1402.5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>344.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>310,-1418.5,323,-1418.5</points>
<connection>
<GID>267</GID>
<name>J</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354,-1401.5,354,-1401</points>
<intersection>-1401.5 2</intersection>
<intersection>-1401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>354,-1401,545,-1401</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>354 0</intersection>
<intersection>545 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>351,-1401.5,354,-1401.5</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>354 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>545,-1401,545,-272.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-1401 1</intersection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333.5,-1424,333.5,-1418.5</points>
<intersection>-1424 2</intersection>
<intersection>-1418.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>329,-1418.5,333.5,-1418.5</points>
<connection>
<GID>267</GID>
<name>Q</name></connection>
<intersection>333.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>333.5,-1424,338.5,-1424</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>333.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-1576.5,277,-1565</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>-1565 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-1565,354,-1565</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,-1564,363,-1425</points>
<intersection>-1564 2</intersection>
<intersection>-1475.5 3</intersection>
<intersection>-1425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,-1425,363,-1425</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>360,-1564,363,-1564</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>363,-1475.5,391,-1475.5</points>
<intersection>363 0</intersection>
<intersection>391 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>391,-1555.5,391,-1475.5</points>
<intersection>-1555.5 5</intersection>
<intersection>-1545.5 7</intersection>
<intersection>-1536 9</intersection>
<intersection>-1527.5 11</intersection>
<intersection>-1519 13</intersection>
<intersection>-1475.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>372,-1555.5,391,-1555.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>391 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>373.5,-1545.5,391,-1545.5</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<intersection>391 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>374,-1536,391,-1536</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>391 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>373.5,-1527.5,391,-1527.5</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>391 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>373,-1519,391,-1519</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<intersection>391 4</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-1576.5,290.5,-1556.5</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>-1556.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-1556.5,366,-1556.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-1576.5,303.5,-1546.5</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>-1546.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-1546.5,367.5,-1546.5</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-1576.5,316.5,-1537</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>-1537 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316.5,-1537,368,-1537</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,-1577,329,-1528.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>-1528.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>329,-1528.5,367.5,-1528.5</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<intersection>329 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-1577,341.5,-1520</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>-1520 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>341.5,-1520,367,-1520</points>
<connection>
<GID>477</GID>
<name>OUT</name></connection>
<intersection>341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-1628.5,350,-1628</points>
<intersection>-1628.5 1</intersection>
<intersection>-1628 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347.5,-1628.5,350,-1628.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>350,-1628,353,-1628</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>178,-658.5,237,-658.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<connection>
<GID>222</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>319,-1637.5,560.5,-1637.5</points>
<connection>
<GID>636</GID>
<name>OUT</name></connection>
<intersection>351 5</intersection>
<intersection>560.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>560.5,-1637.5,560.5,188.5</points>
<intersection>-1637.5 1</intersection>
<intersection>-273 9</intersection>
<intersection>188.5 7</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>351,-1637.5,351,-1630</points>
<intersection>-1637.5 1</intersection>
<intersection>-1630 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>351,-1630,353,-1630</points>
<connection>
<GID>544</GID>
<name>IN_1</name></connection>
<intersection>351 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-244,188.5,560.5,188.5</points>
<intersection>-244 8</intersection>
<intersection>560.5 2</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-244,174,-244,188.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>188.5 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>559,-273,560.5,-273</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>560.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-1629,557,-1629</points>
<connection>
<GID>544</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>557 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>557,-1629,557,-273</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>-1629 1</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519,-266.5,519,-260</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>-260 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>535,-260,535,-254</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>-260 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>519,-260,535,-260</points>
<intersection>519 0</intersection>
<intersection>535 1</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,-266.5,533,-261</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>-261 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>537,-261,537,-254</points>
<connection>
<GID>604</GID>
<name>IN_1</name></connection>
<intersection>-261 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>533,-261,537,-261</points>
<intersection>533 0</intersection>
<intersection>537 1</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-266.5,546,-260</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>-260 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>539,-260,539,-254</points>
<connection>
<GID>604</GID>
<name>IN_2</name></connection>
<intersection>-260 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>539,-260,546,-260</points>
<intersection>539 1</intersection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>558,-267,558,-258</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<intersection>-258 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>541,-258,541,-254</points>
<connection>
<GID>604</GID>
<name>IN_3</name></connection>
<intersection>-258 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>541,-258,558,-258</points>
<intersection>541 1</intersection>
<intersection>558 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>473,-249.5,473,-240.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>-240.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>499,-240.5,499,-232</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>-240.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>473,-240.5,499,-240.5</points>
<intersection>473 0</intersection>
<intersection>499 1</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,-240,501,-232</points>
<connection>
<GID>644</GID>
<name>IN_1</name></connection>
<intersection>-240 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>538,-248,538,-240</points>
<connection>
<GID>604</GID>
<name>OUT</name></connection>
<intersection>-240 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>501,-240,538,-240</points>
<intersection>501 0</intersection>
<intersection>538 1</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-694.5,260,-658.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>-658.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-658.5,260,-658.5</points>
<connection>
<GID>222</GID>
<name>Q</name></connection>
<intersection>260 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177.5,-648.5,224,-648.5</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<connection>
<GID>223</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,-694.5,273.5,-648.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>-648.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,-648.5,273.5,-648.5</points>
<connection>
<GID>223</GID>
<name>Q</name></connection>
<intersection>273.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>176,-637.5,211,-637.5</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<connection>
<GID>224</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-694.5,286.5,-637.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>-637.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,-637.5,286.5,-637.5</points>
<connection>
<GID>224</GID>
<name>Q</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175.5,-628.5,203.5,-628.5</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<connection>
<GID>226</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299.5,-694.5,299.5,-628.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-628.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209.5,-628.5,299.5,-628.5</points>
<connection>
<GID>226</GID>
<name>Q</name></connection>
<intersection>299.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,-621,195,-621</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<connection>
<GID>227</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-695,312,-621</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>-621 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,-621,312,-621</points>
<connection>
<GID>227</GID>
<name>Q</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,-613.5,186,-613.5</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<connection>
<GID>228</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,-695,324.5,-613.5</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>-613.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-613.5,324.5,-613.5</points>
<connection>
<GID>228</GID>
<name>Q</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-660.5,180.5,-609.5</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>-660.5 7</intersection>
<intersection>-650.5 5</intersection>
<intersection>-639.5 8</intersection>
<intersection>-630.5 3</intersection>
<intersection>-623 9</intersection>
<intersection>-615.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,-615.5,186,-615.5</points>
<connection>
<GID>228</GID>
<name>clock</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>180.5,-630.5,203.5,-630.5</points>
<connection>
<GID>226</GID>
<name>clock</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>180.5,-650.5,224,-650.5</points>
<connection>
<GID>223</GID>
<name>clock</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>180.5,-660.5,237,-660.5</points>
<connection>
<GID>222</GID>
<name>clock</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>180.5,-639.5,211,-639.5</points>
<connection>
<GID>224</GID>
<name>clock</name></connection>
<intersection>180.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>180.5,-623,195,-623</points>
<connection>
<GID>227</GID>
<name>clock</name></connection>
<intersection>180.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,-67,502,91.5</points>
<intersection>-67 2</intersection>
<intersection>91.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>500,-226,500,-67</points>
<connection>
<GID>644</GID>
<name>OUT</name></connection>
<intersection>-67 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>500,-67,502,-67</points>
<intersection>500 1</intersection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>22,91.5,502,91.5</points>
<connection>
<GID>431</GID>
<name>clear</name></connection>
<intersection>502 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-946.5,152,-793</points>
<intersection>-946.5 13</intersection>
<intersection>-856.5 1</intersection>
<intersection>-846.5 3</intersection>
<intersection>-835.5 5</intersection>
<intersection>-826.5 7</intersection>
<intersection>-819 9</intersection>
<intersection>-793 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,-856.5,182.5,-856.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>152,-846.5,182,-846.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>152,-835.5,180.5,-835.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>152,-826.5,180,-826.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-819,179,-819</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>152,-793,316,-793</points>
<intersection>152 0</intersection>
<intersection>152.5 17</intersection>
<intersection>178 16</intersection>
<intersection>316 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>152,-946.5,335.5,-946.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>152 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>316,-793,316,-775</points>
<intersection>-793 11</intersection>
<intersection>-775 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>316,-775,325.5,-775</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>316 14</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>178,-811.5,178,-793</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>-793 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>152.5,-793,152.5,-788</points>
<connection>
<GID>1833</GID>
<name>OUT</name></connection>
<intersection>-793 11</intersection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-903,271.5,-899.5</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>-903 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271.5,-903,272.5,-903</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285,-903.5,285,-899.5</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>285,-903.5,288.5,-903.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>285 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298,-903.5,298,-899.5</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>298,-903.5,302,-903.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>298 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-903.5,314,-899.5</points>
<intersection>-903.5 1</intersection>
<intersection>-899.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-903.5,317,-903.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>311,-899.5,314,-899.5</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323.5,-902,323.5,-900</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>-902 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,-902,327.5,-902</points>
<intersection>323.5 0</intersection>
<intersection>327.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>327.5,-903.5,327.5,-902</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>-902 1</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336,-902,336,-900</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>-902 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336,-902,340.5,-902</points>
<intersection>336 0</intersection>
<intersection>340.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>340.5,-903.5,340.5,-902</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>-902 1</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-911,282.5,-903</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>-903 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278.5,-903,282.5,-903</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-911,297.5,-903.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,-903.5,297.5,-903.5</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-911,312.5,-903.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308,-903.5,312.5,-903.5</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324,-910.5,324,-903.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,-903.5,324,-903.5</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>324 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-911,337,-903.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>333.5,-903.5,337,-903.5</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>337 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-910.5,350,-903.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>-903.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>346.5,-903.5,350,-903.5</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-920.5,282.5,-915</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>-920.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>297.5,-926.5,297.5,-920.5</points>
<connection>
<GID>291</GID>
<name>IN_3</name></connection>
<intersection>-920.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>282.5,-920.5,297.5,-920.5</points>
<intersection>282.5 0</intersection>
<intersection>297.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-920,297.5,-915</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>-920 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>299.5,-926.5,299.5,-920</points>
<connection>
<GID>291</GID>
<name>IN_2</name></connection>
<intersection>-920 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>297.5,-920,299.5,-920</points>
<intersection>297.5 0</intersection>
<intersection>299.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-920.5,312.5,-915</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>-920.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>301.5,-926.5,301.5,-920.5</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>-920.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-920.5,312.5,-920.5</points>
<intersection>301.5 1</intersection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324,-921.5,324,-914.5</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>-921.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>303.5,-926.5,303.5,-921.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>-921.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-921.5,324,-921.5</points>
<intersection>303.5 1</intersection>
<intersection>324 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-920,337,-915</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-920 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>336,-925.5,336,-920</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>-920 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>336,-920,337,-920</points>
<intersection>336 1</intersection>
<intersection>337 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-920,350,-914.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>-920 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>338,-925.5,338,-920</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-920 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>338,-920,350,-920</points>
<intersection>338 1</intersection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300.5,-935.5,300.5,-932.5</points>
<connection>
<GID>291</GID>
<name>OUT</name></connection>
<intersection>-935.5 2</intersection>
<intersection>-935 8</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>313.5,-948.5,313.5,-935.5</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>-943.5 7</intersection>
<intersection>-935.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-935.5,313.5,-935.5</points>
<intersection>300.5 0</intersection>
<intersection>313.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>313.5,-943.5,325,-943.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>313.5 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>245,-935,300.5,-935</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>300.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-935,337,-931.5</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>-935 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>315.5,-948.5,315.5,-935</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>-945.5 6</intersection>
<intersection>-939.5 7</intersection>
<intersection>-935 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>315.5,-935,337,-935</points>
<intersection>315.5 1</intersection>
<intersection>337 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>315.5,-945.5,325,-945.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>315.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>204.5,-939.5,315.5,-939.5</points>
<intersection>204.5 8</intersection>
<intersection>315.5 1</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>204.5,-939.5,204.5,-937</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-939.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,-857.5,247.5,-857.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<connection>
<GID>305</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-893.5,270.5,-857.5</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>-857.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253.5,-857.5,270.5,-857.5</points>
<connection>
<GID>305</GID>
<name>Q</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188,-847.5,234.5,-847.5</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-893.5,284,-847.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>-847.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240.5,-847.5,284,-847.5</points>
<connection>
<GID>306</GID>
<name>Q</name></connection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186.5,-836.5,221.5,-836.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<connection>
<GID>307</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297,-893.5,297,-836.5</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>-836.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,-836.5,297,-836.5</points>
<connection>
<GID>307</GID>
<name>Q</name></connection>
<intersection>297 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>186,-827.5,214,-827.5</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<connection>
<GID>309</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-893.5,310,-827.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>-827.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-827.5,310,-827.5</points>
<connection>
<GID>309</GID>
<name>Q</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-820,205.5,-820</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<connection>
<GID>310</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322.5,-894,322.5,-820</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>-820 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-820,322.5,-820</points>
<connection>
<GID>310</GID>
<name>Q</name></connection>
<intersection>322.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184,-812.5,196.5,-812.5</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<connection>
<GID>311</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-894,335,-812.5</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>-812.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-812.5,335,-812.5</points>
<connection>
<GID>311</GID>
<name>Q</name></connection>
<intersection>335 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-859.5,191.5,-808.5</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>-859.5 7</intersection>
<intersection>-849.5 5</intersection>
<intersection>-838.5 8</intersection>
<intersection>-829.5 3</intersection>
<intersection>-822 9</intersection>
<intersection>-814.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-814.5,196.5,-814.5</points>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191.5,-829.5,214,-829.5</points>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>191.5,-849.5,234.5,-849.5</points>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>191.5,-859.5,247.5,-859.5</points>
<connection>
<GID>305</GID>
<name>clock</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>191.5,-838.5,221.5,-838.5</points>
<connection>
<GID>307</GID>
<name>clock</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>191.5,-822,205.5,-822</points>
<connection>
<GID>310</GID>
<name>clock</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,-377,308.5,-372</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>-377 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>307.5,-382.5,307.5,-377</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>-377 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-377,308.5,-377</points>
<intersection>307.5 1</intersection>
<intersection>308.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,-377,321.5,-371.5</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>-377 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>309.5,-382.5,309.5,-377</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-377 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-377,321.5,-377</points>
<intersection>309.5 1</intersection>
<intersection>321.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-392.5,272,-389.5</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>-392.5 2</intersection>
<intersection>-389.5 5</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>286.5,-400.5,286.5,-392.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>-394.5 3</intersection>
<intersection>-392.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>272,-392.5,286.5,-392.5</points>
<intersection>272 0</intersection>
<intersection>286.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286.5,-394.5,325,-394.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>286.5 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>252,-389.5,272,-389.5</points>
<intersection>252 6</intersection>
<intersection>272 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>252,-390,252,-389.5</points>
<intersection>-390 10</intersection>
<intersection>-389.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>164,-390,252,-390</points>
<connection>
<GID>1801</GID>
<name>IN_0</name></connection>
<intersection>252 6</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,-392.5,308.5,-388.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>-392.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>288.5,-400.5,288.5,-392.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>-395.5 4</intersection>
<intersection>-392.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>288.5,-392.5,325,-392.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>288.5 1</intersection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>154,-395.5,288.5,-395.5</points>
<intersection>154 5</intersection>
<intersection>288.5 1</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>154,-395.5,154,-391</points>
<intersection>-395.5 4</intersection>
<intersection>-391 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>152,-391,154,-391</points>
<connection>
<GID>1797</GID>
<name>IN_0</name></connection>
<intersection>154 5</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-1168.5,146,-1005.5</points>
<connection>
<GID>1837</GID>
<name>OUT</name></connection>
<intersection>-1168.5 13</intersection>
<intersection>-1078.5 1</intersection>
<intersection>-1068.5 3</intersection>
<intersection>-1057.5 5</intersection>
<intersection>-1048.5 7</intersection>
<intersection>-1041 9</intersection>
<intersection>-1009 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146,-1078.5,176,-1078.5</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>146,-1068.5,175.5,-1068.5</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>146,-1057.5,174,-1057.5</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>146,-1048.5,173.5,-1048.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>146,-1041,172.5,-1041</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>146,-1009,338.5,-1009</points>
<intersection>146 0</intersection>
<intersection>171.5 15</intersection>
<intersection>338.5 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>146,-1168.5,331,-1168.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>146 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>338.5,-1009,338.5,-970.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>-1009 11</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>171.5,-1033.5,171.5,-1009</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>-1009 11</intersection></vsegment></shape></wire>
<wire>
<ID>1835</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,-347,337.5,-297.5</points>
<intersection>-347 1</intersection>
<intersection>-315 3</intersection>
<intersection>-297.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>334.5,-347,337.5,-347</points>
<connection>
<GID>2094</GID>
<name>IN_1</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>335.5,-297.5,337.5,-297.5</points>
<connection>
<GID>2092</GID>
<name>OUT</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>337.5,-315,361,-315</points>
<intersection>337.5 0</intersection>
<intersection>349 12</intersection>
<intersection>361 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>361,-344,361,-315</points>
<intersection>-344 7</intersection>
<intersection>-336.5 6</intersection>
<intersection>-328.5 9</intersection>
<intersection>-322.5 11</intersection>
<intersection>-315 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>347.5,-336.5,361,-336.5</points>
<connection>
<GID>2098</GID>
<name>IN_1</name></connection>
<intersection>361 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>348,-344,361,-344</points>
<connection>
<GID>2096</GID>
<name>IN_1</name></connection>
<intersection>361 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>348.5,-328.5,361,-328.5</points>
<connection>
<GID>2100</GID>
<name>IN_1</name></connection>
<intersection>361 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>348.5,-322.5,361,-322.5</points>
<connection>
<GID>2102</GID>
<name>IN_1</name></connection>
<intersection>361 4</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>349,-317,349,-315</points>
<connection>
<GID>2104</GID>
<name>IN_1</name></connection>
<intersection>-315 3</intersection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265,-1125,265,-1121.5</points>
<connection>
<GID>534</GID>
<name>OUT</name></connection>
<intersection>-1125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265,-1125,266,-1125</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>265 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-1125.5,278.5,-1121.5</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278.5,-1125.5,282,-1125.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1836</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-350.5,244,-348</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>-348 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-348,328.5,-348</points>
<connection>
<GID>2094</GID>
<name>OUT</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>1837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-350.5,257.5,-345</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-345 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-345,342,-345</points>
<connection>
<GID>2096</GID>
<name>OUT</name></connection>
<intersection>257.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-350.5,270.5,-337.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>-337.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-337.5,341.5,-337.5</points>
<connection>
<GID>2098</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-1125.5,291.5,-1121.5</points>
<connection>
<GID>538</GID>
<name>OUT</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,-1125.5,296,-1125.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,-350.5,283.5,-329.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>-329.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283.5,-329.5,342.5,-329.5</points>
<connection>
<GID>2100</GID>
<name>OUT</name></connection>
<intersection>283.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-1125.5,307.5,-1121.5</points>
<intersection>-1125.5 1</intersection>
<intersection>-1121.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>307.5,-1125.5,310.5,-1125.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>307.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>304.5,-1121.5,307.5,-1121.5</points>
<connection>
<GID>539</GID>
<name>OUT</name></connection>
<intersection>307.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-351,296,-323.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>-323.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>296,-323.5,342.5,-323.5</points>
<connection>
<GID>2102</GID>
<name>OUT</name></connection>
<intersection>296 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-1124,317,-1122</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<intersection>-1124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-1124,321,-1124</points>
<intersection>317 0</intersection>
<intersection>321 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>321,-1125.5,321,-1124</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-1124 1</intersection></vsegment></shape></wire>
<wire>
<ID>1841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,-351,308.5,-318</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>-318 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308.5,-318,343,-318</points>
<connection>
<GID>2104</GID>
<name>OUT</name></connection>
<intersection>308.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-188.5,123.5,-139</points>
<connection>
<GID>1818</GID>
<name>OUT</name></connection>
<intersection>-188.5 1</intersection>
<intersection>-178.5 3</intersection>
<intersection>-167.5 5</intersection>
<intersection>-158.5 7</intersection>
<intersection>-151 9</intersection>
<intersection>-143.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-188.5,154.5,-188.5</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection>
<intersection>139 12</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123.5,-178.5,154,-178.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>123.5,-167.5,152.5,-167.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>123.5,-158.5,152,-158.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>123.5,-151,151,-151</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>123.5,-143.5,150,-143.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>139,-284.5,139,-188.5</points>
<intersection>-284.5 13</intersection>
<intersection>-188.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>139,-284.5,320,-284.5</points>
<intersection>139 12</intersection>
<intersection>320 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>320,-284.5,320,-284</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>-284.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>1842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347.5,-400.5,347.5,-400</points>
<intersection>-400.5 2</intersection>
<intersection>-400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345,-400,347.5,-400</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>347.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347.5,-400.5,350.5,-400.5</points>
<connection>
<GID>2106</GID>
<name>IN_0</name></connection>
<intersection>347.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-1124,329.5,-1122</points>
<connection>
<GID>542</GID>
<name>OUT</name></connection>
<intersection>-1124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>329.5,-1124,334,-1124</points>
<intersection>329.5 0</intersection>
<intersection>334 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>334,-1125.5,334,-1124</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>-1124 1</intersection></vsegment></shape></wire>
<wire>
<ID>1843</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>287.5,-406.5,469,-406.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>302 6</intersection>
<intersection>350.5 5</intersection>
<intersection>469 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>469,-406.5,469,-271.5</points>
<connection>
<GID>2108</GID>
<name>IN_1</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>350.5,-406.5,350.5,-402.5</points>
<connection>
<GID>2106</GID>
<name>IN_1</name></connection>
<intersection>-406.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>302,-408,302,-406.5</points>
<connection>
<GID>7</GID>
<name>J</name></connection>
<intersection>-406.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-1133,276,-1125</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-1125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,-1125,276,-1125</points>
<connection>
<GID>578</GID>
<name>OUT_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>1844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360.5,-401.5,360.5,-400</points>
<intersection>-401.5 2</intersection>
<intersection>-400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360.5,-400,467,-400</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>360.5 0</intersection>
<intersection>467 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>356.5,-401.5,360.5,-401.5</points>
<connection>
<GID>2106</GID>
<name>OUT</name></connection>
<intersection>360.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>467,-400,467,-271.5</points>
<connection>
<GID>2108</GID>
<name>IN_0</name></connection>
<intersection>-400 1</intersection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243.5,-235,243.5,-231.5</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243.5,-235,244.5,-235</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>243.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-235.5,257,-231.5</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-235.5,260.5,-235.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-235.5,270,-231.5</points>
<connection>
<GID>516</GID>
<name>OUT</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-235.5,274,-235.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-235.5,286,-231.5</points>
<intersection>-235.5 1</intersection>
<intersection>-231.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-235.5,289,-235.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>283,-231.5,286,-231.5</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<intersection>286 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-234,295.5,-232</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>-234 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-234,299.5,-234</points>
<intersection>295.5 0</intersection>
<intersection>299.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>299.5,-235.5,299.5,-234</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>-234 1</intersection></vsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-234,308,-232</points>
<connection>
<GID>521</GID>
<name>OUT</name></connection>
<intersection>-234 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308,-234,312.5,-234</points>
<intersection>308 0</intersection>
<intersection>312.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>312.5,-235.5,312.5,-234</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>-234 1</intersection></vsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254.5,-243,254.5,-235</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>-235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-235,254.5,-235</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<intersection>254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-243,269.5,-235.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266.5,-235.5,269.5,-235.5</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-243,284.5,-235.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280,-235.5,284.5,-235.5</points>
<connection>
<GID>403</GID>
<name>OUT_0</name></connection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-242.5,296,-235.5</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295,-235.5,296,-235.5</points>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection>
<intersection>296 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-243,309,-235.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>305.5,-235.5,309,-235.5</points>
<connection>
<GID>415</GID>
<name>OUT_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,-242.5,322,-235.5</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-235.5,322,-235.5</points>
<connection>
<GID>422</GID>
<name>OUT_0</name></connection>
<intersection>322 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254.5,-252.5,254.5,-247</points>
<connection>
<GID>427</GID>
<name>OUT_0</name></connection>
<intersection>-252.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>269.5,-258.5,269.5,-252.5</points>
<connection>
<GID>456</GID>
<name>IN_3</name></connection>
<intersection>-252.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>254.5,-252.5,269.5,-252.5</points>
<intersection>254.5 0</intersection>
<intersection>269.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-252,269.5,-247</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<intersection>-252 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>271.5,-258.5,271.5,-252</points>
<connection>
<GID>456</GID>
<name>IN_2</name></connection>
<intersection>-252 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-252,271.5,-252</points>
<intersection>269.5 0</intersection>
<intersection>271.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-252.5,284.5,-247</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<intersection>-252.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>273.5,-258.5,273.5,-252.5</points>
<connection>
<GID>456</GID>
<name>IN_1</name></connection>
<intersection>-252.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>273.5,-252.5,284.5,-252.5</points>
<intersection>273.5 1</intersection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-253.5,296,-246.5</points>
<connection>
<GID>435</GID>
<name>OUT_0</name></connection>
<intersection>-253.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>275.5,-258.5,275.5,-253.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>-253.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>275.5,-253.5,296,-253.5</points>
<intersection>275.5 1</intersection>
<intersection>296 0</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-252,309,-247</points>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection>
<intersection>-252 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>308,-257.5,308,-252</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<intersection>-252 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308,-252,309,-252</points>
<intersection>308 1</intersection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,-252,322,-246.5</points>
<connection>
<GID>440</GID>
<name>OUT_0</name></connection>
<intersection>-252 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>310,-257.5,310,-252</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>-252 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>310,-252,322,-252</points>
<intersection>310 1</intersection>
<intersection>322 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-268,272.5,-264.5</points>
<connection>
<GID>456</GID>
<name>OUT</name></connection>
<intersection>-268 9</intersection>
<intersection>-267.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>285.5,-280.5,285.5,-267.5</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>-275.5 7</intersection>
<intersection>-267.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>272.5,-267.5,285.5,-267.5</points>
<intersection>272.5 0</intersection>
<intersection>285.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>285.5,-275.5,297,-275.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>285.5 1</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>175.5,-268,272.5,-268</points>
<connection>
<GID>1795</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-267,309,-263.5</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>-267 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>287.5,-280.5,287.5,-267</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>-277.5 6</intersection>
<intersection>-272 7</intersection>
<intersection>-267 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>287.5,-267,309,-267</points>
<intersection>287.5 1</intersection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>287.5,-277.5,297,-277.5</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>287.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>164.5,-272,287.5,-272</points>
<connection>
<GID>1785</GID>
<name>IN_0</name></connection>
<intersection>287.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-1133,291,-1125.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,-1125.5,291,-1125.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306,-1133,306,-1125.5</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,-1125.5,306,-1125.5</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>306 0</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-1132.5,317.5,-1125.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316.5,-1125.5,317.5,-1125.5</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-311.5,-6.5,-304,-6.5</points>
<connection>
<GID>512</GID>
<name>OUT_0</name></connection>
<connection>
<GID>511</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-262,-8.5,-254,-8.5</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<connection>
<GID>523</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-258,-17,-258,-11.5</points>
<intersection>-17 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-258,-11.5,-254,-11.5</points>
<connection>
<GID>523</GID>
<name>clock</name></connection>
<intersection>-258 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-304,-17,-258,-17</points>
<intersection>-304 3</intersection>
<intersection>-262 4</intersection>
<intersection>-258 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-304,-17,-304,-9.5</points>
<connection>
<GID>511</GID>
<name>clock</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-262,-17,-262,-14</points>
<connection>
<GID>524</GID>
<name>CLK</name></connection>
<intersection>-17 2</intersection></vsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-283.5,-20.5,-283.5,-0.5</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-283.5,-20.5,-248,-20.5</points>
<intersection>-283.5 0</intersection>
<intersection>-248 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-248,-20.5,-248,-11.5</points>
<connection>
<GID>523</GID>
<name>OUTINV_0</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-285.5,-6.5,-285.5,-0.5</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-298,-6.5,-285.5,-6.5</points>
<connection>
<GID>511</GID>
<name>OUT_0</name></connection>
<intersection>-285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-284.5,5.5,-284.5,157.5</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<intersection>157.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-284.5,157.5,-248,157.5</points>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<intersection>-284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-298,-9.5,-292.5,-9.5</points>
<connection>
<GID>511</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>520</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-251,-49.5,-251,-14.5</points>
<connection>
<GID>523</GID>
<name>clear</name></connection>
<intersection>-49.5 3</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-288.5,-22,-251,-22</points>
<intersection>-288.5 2</intersection>
<intersection>-251 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-288.5,-22,-288.5,-9.5</points>
<connection>
<GID>520</GID>
<name>OUT_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-251,-49.5,-235.5,-49.5</points>
<connection>
<GID>388</GID>
<name>clear</name></connection>
<intersection>-251 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-67,53,-11.5</points>
<intersection>-67 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-11.5,53,-11.5</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-172,-67,53,-67</points>
<intersection>-172 15</intersection>
<intersection>-122.5 14</intersection>
<intersection>-96.5 10</intersection>
<intersection>-66.5 18</intersection>
<intersection>-28 16</intersection>
<intersection>20.5 17</intersection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-96.5,-67,-96.5,-41</points>
<connection>
<GID>359</GID>
<name>clear</name></connection>
<intersection>-67 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-122.5,-67,-122.5,-41.5</points>
<connection>
<GID>357</GID>
<name>clear</name></connection>
<intersection>-67 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-172,-67,-172,-41</points>
<connection>
<GID>355</GID>
<name>clear</name></connection>
<intersection>-67 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-28,-67,-28,-43.5</points>
<connection>
<GID>363</GID>
<name>clear</name></connection>
<intersection>-67 2</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>20.5,-67,20.5,-44</points>
<connection>
<GID>365</GID>
<name>clear</name></connection>
<intersection>-67 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-66.5,-67,-66.5,-41.5</points>
<connection>
<GID>361</GID>
<name>clear</name></connection>
<intersection>-67 2</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-163,-79.5,-163,-29</points>
<intersection>-79.5 8</intersection>
<intersection>-73.5 5</intersection>
<intersection>-64 3</intersection>
<intersection>-35 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-163,-29,-158.5,-29</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>-163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-169,-35,-163,-35</points>
<connection>
<GID>355</GID>
<name>Q</name></connection>
<intersection>-163 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-163,-64,40,-64</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-163 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-163,-73.5,-144,-73.5</points>
<intersection>-163 0</intersection>
<intersection>-144 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-144,-106,-144,-73.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>-73.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-163,-79.5,-157,-79.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-163 0</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-167,-44.5,-167,-39</points>
<intersection>-44.5 3</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-169,-39,-167,-39</points>
<connection>
<GID>355</GID>
<name>nQ</name></connection>
<intersection>-167 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-167,-44.5,-159.5,-44.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>-167 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148.5,-36.5,-148.5,-27</points>
<intersection>-36.5 1</intersection>
<intersection>-28 2</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-148.5,-36.5,-144.5,-36.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>-148.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-152.5,-28,-148.5,-28</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<intersection>-148.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-148.5,-27,-117.5,-27</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>-148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148,-47.5,-148,-38.5</points>
<intersection>-47.5 2</intersection>
<intersection>-45.5 3</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-148,-38.5,-144.5,-38.5</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<intersection>-148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-148,-47.5,-115,-47.5</points>
<connection>
<GID>371</GID>
<name>IN_1</name></connection>
<intersection>-148 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-153.5,-45.5,-148,-45.5</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<intersection>-148 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-118.5,-105.5,-118.5,-29</points>
<intersection>-105.5 9</intersection>
<intersection>-79 5</intersection>
<intersection>-63 3</intersection>
<intersection>-35.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-118.5,-29,-117.5,-29</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>-118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-119.5,-35.5,-118.5,-35.5</points>
<connection>
<GID>357</GID>
<name>Q</name></connection>
<intersection>-118.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-118.5,-63,40,-63</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>-118.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118.5,-79,-114,-79</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>-118.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-131.5,-105.5,-118.5,-105.5</points>
<intersection>-131.5 10</intersection>
<intersection>-118.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-131.5,-107,-131.5,-105.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>-105.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148,-347,-148,-79.5</points>
<intersection>-347 12</intersection>
<intersection>-191 5</intersection>
<intersection>-94.5 10</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-151,-79.5,-148,-79.5</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>-148 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-148,-191,154.5,-191</points>
<intersection>-148 0</intersection>
<intersection>154.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>154.5,-191,154.5,-190.5</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>-191 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-148,-94.5,59.5,-94.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-148 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-148,-347,151.5,-347</points>
<connection>
<GID>528</GID>
<name>IN_1</name></connection>
<intersection>-148 0</intersection>
<intersection>-147.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-147.5,-858.5,-147.5,-347</points>
<intersection>-858.5 19</intersection>
<intersection>-659.5 17</intersection>
<intersection>-477.5 15</intersection>
<intersection>-347 12</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-147.5,-477.5,164,-477.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>-147.5 14</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-147.5,-659.5,172,-659.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>-147.5 14</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-147.5,-858.5,182.5,-858.5</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-147.5 14</intersection>
<intersection>-146.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-146.5,-1080.5,-146.5,-858.5</points>
<intersection>-1080.5 21</intersection>
<intersection>-858.5 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-146.5,-1080.5,176,-1080.5</points>
<connection>
<GID>571</GID>
<name>IN_1</name></connection>
<intersection>-146.5 20</intersection>
<intersection>-145.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-145.5,-1314.5,-145.5,-1080.5</points>
<intersection>-1314.5 23</intersection>
<intersection>-1080.5 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>-145.5,-1314.5,178,-1314.5</points>
<connection>
<GID>614</GID>
<name>IN_1</name></connection>
<intersection>-145.5 22</intersection>
<intersection>-144 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-144,-1541.5,-144,-1314.5</points>
<intersection>-1541.5 25</intersection>
<intersection>-1314.5 23</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>-144,-1541.5,187,-1541.5</points>
<connection>
<GID>656</GID>
<name>IN_1</name></connection>
<intersection>-144 24</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110,-28.5,-110,-28</points>
<intersection>-28.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111.5,-28,-110,-28</points>
<connection>
<GID>370</GID>
<name>OUT</name></connection>
<intersection>-110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-110,-28.5,-88,-28.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>-110 0</intersection>
<intersection>-108 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-108,-35.5,-108,-28.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-28.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-117,-45.5,-117,-39.5</points>
<intersection>-45.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-119.5,-39.5,-117,-39.5</points>
<connection>
<GID>357</GID>
<name>nQ</name></connection>
<intersection>-117 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-117,-45.5,-115,-45.5</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-117 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108.5,-49,-108.5,-37.5</points>
<intersection>-49 3</intersection>
<intersection>-46.5 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109,-46.5,-108.5,-46.5</points>
<connection>
<GID>371</GID>
<name>OUT</name></connection>
<intersection>-108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-108.5,-37.5,-108,-37.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>-108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108.5,-49,-85.5,-49</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<intersection>-108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91.5,-106,-91.5,-8.5</points>
<intersection>-106 13</intersection>
<intersection>-79 9</intersection>
<intersection>-62 2</intersection>
<intersection>-35 1</intersection>
<intersection>-30.5 5</intersection>
<intersection>-8.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-35,-91.5,-35</points>
<connection>
<GID>359</GID>
<name>Q</name></connection>
<intersection>-91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-91.5,-62,40,-62</points>
<connection>
<GID>387</GID>
<name>IN_2</name></connection>
<intersection>-91.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-91.5,-30.5,-88,-30.5</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>-91.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-91.5,-8.5,42,-8.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-91.5,-79,-84.5,-79</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>-91.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-91.5,-106,-67.5,-106</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>-91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,-29.5,-61.5,-29.5</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-79.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-79.5,-36,-79.5,-29.5</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79.5,-49,-79.5,-38</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-79.5,-49,-60,-49</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>-79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90,-47,-90,-39</points>
<intersection>-47 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-39,-90,-39</points>
<connection>
<GID>359</GID>
<name>nQ</name></connection>
<intersection>-90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90,-47,-85.5,-47</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-90 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-79,-63.5,-10.5</points>
<connection>
<GID>361</GID>
<name>Q</name></connection>
<intersection>-79 10</intersection>
<intersection>-61 2</intersection>
<intersection>-31.5 6</intersection>
<intersection>-10.5 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-63.5,-61,40,-61</points>
<connection>
<GID>387</GID>
<name>IN_3</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-63.5,-31.5,-61.5,-31.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-63.5,-10.5,42,-10.5</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-63.5,-79,-56,-79</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-63.5 0</intersection>
<intersection>-60.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-60.5,-106,-60.5,-79</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>-79 10</intersection></vsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-47,-62.5,-39.5</points>
<intersection>-47 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-39.5,-62.5,-39.5</points>
<connection>
<GID>361</GID>
<name>nQ</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62.5,-47,-60,-47</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-36.5,-52.5,-28.5</points>
<intersection>-36.5 2</intersection>
<intersection>-30.5 1</intersection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,-30.5,-52.5,-30.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-36.5,-50.5,-36.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-52.5,-28.5,-14.5,-28.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-48,-52,-38.5</points>
<intersection>-48 1</intersection>
<intersection>-38.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-48,-14,-48</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-52,-38.5,-50.5,-38.5</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-105.5,-20,-12.5</points>
<intersection>-105.5 14</intersection>
<intersection>-79 9</intersection>
<intersection>-60 3</intersection>
<intersection>-37.5 1</intersection>
<intersection>-30.5 10</intersection>
<intersection>-12.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-37.5,-20,-37.5</points>
<connection>
<GID>363</GID>
<name>Q</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-20,-60,40,-60</points>
<connection>
<GID>387</GID>
<name>IN_4</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-20,-12.5,42,-12.5</points>
<connection>
<GID>352</GID>
<name>IN_2</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-20,-79,-10,-79</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-20,-30.5,-14.5,-30.5</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-20,-105.5,-3,-105.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-46,-22.5,-41.5</points>
<intersection>-46 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-41.5,-22.5,-41.5</points>
<connection>
<GID>363</GID>
<name>nQ</name></connection>
<intersection>-22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,-46,-14,-46</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-37,-7.5,-29.5</points>
<intersection>-37 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-29.5,-7.5,-29.5</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-37,-6.5,-37</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-47,-7.5,-39</points>
<intersection>-47 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-47,-7.5,-47</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-39,-6.5,-39</points>
<connection>
<GID>385</GID>
<name>IN_1</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-200.5,-56.5,17.5,-56.5</points>
<intersection>-200.5 16</intersection>
<intersection>-183 13</intersection>
<intersection>-126 12</intersection>
<intersection>-100.5 6</intersection>
<intersection>-72.5 7</intersection>
<intersection>-34.5 11</intersection>
<intersection>17.5 28</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-100.5,-56.5,-100.5,-37</points>
<intersection>-56.5 1</intersection>
<intersection>-37 19</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-72.5,-56.5,-72.5,-37.5</points>
<intersection>-56.5 1</intersection>
<intersection>-37.5 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-34.5,-56.5,-34.5,-39.5</points>
<intersection>-56.5 1</intersection>
<intersection>-39.5 18</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-126,-56.5,-126,-37.5</points>
<intersection>-56.5 1</intersection>
<intersection>-37.5 22</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-183,-56.5,-183,-37</points>
<intersection>-56.5 1</intersection>
<intersection>-37 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-72.5,-37.5,-69.5,-37.5</points>
<connection>
<GID>361</GID>
<name>clock</name></connection>
<intersection>-72.5 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-183,-37,-175,-37</points>
<connection>
<GID>355</GID>
<name>clock</name></connection>
<intersection>-183 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-200.5,-86,-200.5,-56.5</points>
<intersection>-86 17</intersection>
<intersection>-57 37</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-200.5,-86,38,-86</points>
<intersection>-200.5 16</intersection>
<intersection>-157 34</intersection>
<intersection>-114 25</intersection>
<intersection>-84.5 26</intersection>
<intersection>-56 24</intersection>
<intersection>-11 23</intersection>
<intersection>38 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-34.5,-39.5,-31,-39.5</points>
<connection>
<GID>363</GID>
<name>clock</name></connection>
<intersection>-34.5 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-100.5,-37,-99.5,-37</points>
<connection>
<GID>359</GID>
<name>clock</name></connection>
<intersection>-100.5 6</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-126,-37.5,-125.5,-37.5</points>
<connection>
<GID>357</GID>
<name>clock</name></connection>
<intersection>-126 12</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-11,-86,-11,-82</points>
<intersection>-86 17</intersection>
<intersection>-82 36</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-56,-86,-56,-82</points>
<connection>
<GID>378</GID>
<name>clock</name></connection>
<intersection>-86 17</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>-114,-86,-114,-82</points>
<connection>
<GID>358</GID>
<name>clock</name></connection>
<intersection>-86 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-84.5,-86,-84.5,-82</points>
<connection>
<GID>366</GID>
<name>clock</name></connection>
<intersection>-86 17</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>17.5,-56.5,17.5,-40</points>
<connection>
<GID>365</GID>
<name>clock</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-157,-86,-157,-82.5</points>
<connection>
<GID>353</GID>
<name>clock</name></connection>
<intersection>-86 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>38,-86,38,-82.5</points>
<connection>
<GID>386</GID>
<name>clock</name></connection>
<intersection>-86 17</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>-11,-82,-10,-82</points>
<connection>
<GID>381</GID>
<name>clock</name></connection>
<intersection>-11 23</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-241.5,-57,-200.5,-57</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<intersection>-239 38</intersection>
<intersection>-200.5 16</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>-239,-57,-239,-46.5</points>
<intersection>-57 37</intersection>
<intersection>-46.5 39</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-239,-46.5,-238.5,-46.5</points>
<connection>
<GID>388</GID>
<name>clock</name></connection>
<intersection>-239 38</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-105,32.5,-14.5</points>
<intersection>-105 9</intersection>
<intersection>-79.5 13</intersection>
<intersection>-59 2</intersection>
<intersection>-38 11</intersection>
<intersection>-14.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-59,40,-59</points>
<connection>
<GID>387</GID>
<name>IN_5</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>32.5,-14.5,42,-14.5</points>
<connection>
<GID>352</GID>
<name>IN_3</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>2.5,-105,32.5,-105</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>23.5,-38,32.5,-38</points>
<connection>
<GID>365</GID>
<name>Q</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>32.5,-79.5,38,-79.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-106.5,-649.5,-106.5,-79</points>
<intersection>-649.5 20</intersection>
<intersection>-467.5 18</intersection>
<intersection>-338.5 16</intersection>
<intersection>-180.5 11</intersection>
<intersection>-93.5 14</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-108,-79,-106.5,-79</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-106.5,-180.5,154,-180.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-106.5,-93.5,59.5,-93.5</points>
<connection>
<GID>390</GID>
<name>IN_1</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-106.5,-338.5,151,-338.5</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-106.5,-467.5,163.5,-467.5</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-106.5,-649.5,171.5,-649.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>-106.5 3</intersection>
<intersection>-106 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>-106,-848.5,-106,-649.5</points>
<intersection>-848.5 22</intersection>
<intersection>-649.5 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>-108,-848.5,182,-848.5</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>-108 23</intersection>
<intersection>-106 21</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-108,-1531.5,-108,-848.5</points>
<intersection>-1531.5 28</intersection>
<intersection>-1304.5 26</intersection>
<intersection>-1070.5 24</intersection>
<intersection>-848.5 22</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-108,-1070.5,175.5,-1070.5</points>
<connection>
<GID>573</GID>
<name>IN_1</name></connection>
<intersection>-108 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-108,-1304.5,177.5,-1304.5</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<intersection>-108 23</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-108,-1531.5,186.5,-1531.5</points>
<connection>
<GID>657</GID>
<name>IN_1</name></connection>
<intersection>-108 23</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-77,-330,-77,-79</points>
<intersection>-330 14</intersection>
<intersection>-169.5 7</intersection>
<intersection>-92.5 12</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-78.5,-79,-77,-79</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<intersection>-77 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-77,-169.5,152.5,-169.5</points>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<intersection>-77 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-77,-92.5,59.5,-92.5</points>
<connection>
<GID>390</GID>
<name>IN_2</name></connection>
<intersection>-77 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-77,-330,150.5,-330</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>-77 3</intersection>
<intersection>-76.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-76.5,-638.5,-76.5,-330</points>
<intersection>-638.5 18</intersection>
<intersection>-456.5 16</intersection>
<intersection>-330 14</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-76.5,-456.5,162,-456.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>-76.5 15</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-76.5,-638.5,170,-638.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>-76.5 15</intersection>
<intersection>-76 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-76,-837.5,-76,-638.5</points>
<intersection>-837.5 20</intersection>
<intersection>-638.5 18</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-76,-837.5,180.5,-837.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>-76 19</intersection>
<intersection>-75.5 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>-75.5,-1059.5,-75.5,-837.5</points>
<intersection>-1059.5 22</intersection>
<intersection>-837.5 20</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>-76,-1059.5,174,-1059.5</points>
<connection>
<GID>574</GID>
<name>IN_1</name></connection>
<intersection>-76 23</intersection>
<intersection>-75.5 21</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-76,-1520.5,-76,-1059.5</points>
<intersection>-1520.5 26</intersection>
<intersection>-1293.5 24</intersection>
<intersection>-1059.5 22</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-76,-1293.5,176,-1293.5</points>
<connection>
<GID>616</GID>
<name>IN_1</name></connection>
<intersection>-76 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-76,-1520.5,185,-1520.5</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<intersection>-76 23</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-50,-447.5,-50,-79</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<intersection>-447.5 19</intersection>
<intersection>-322 17</intersection>
<intersection>-160.5 7</intersection>
<intersection>-91.5 15</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-50,-160.5,152,-160.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>-50 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-50,-91.5,59.5,-91.5</points>
<connection>
<GID>390</GID>
<name>IN_3</name></connection>
<intersection>-50 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-50,-322,150,-322</points>
<connection>
<GID>531</GID>
<name>IN_1</name></connection>
<intersection>-50 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-50,-447.5,161.5,-447.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>-50 3</intersection>
<intersection>-49.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-49.5,-1050.5,-49.5,-447.5</points>
<intersection>-1050.5 25</intersection>
<intersection>-828.5 23</intersection>
<intersection>-629.5 21</intersection>
<intersection>-447.5 19</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-49.5,-629.5,169.5,-629.5</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>-49.5 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-49.5,-828.5,180,-828.5</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>-49.5 20</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-49.5,-1050.5,173.5,-1050.5</points>
<connection>
<GID>575</GID>
<name>IN_1</name></connection>
<intersection>-49.5 20</intersection>
<intersection>-49 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>-49,-1284.5,-49,-1050.5</points>
<intersection>-1284.5 27</intersection>
<intersection>-1050.5 25</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-49.5,-1284.5,175.5,-1284.5</points>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>-49.5 28</intersection>
<intersection>-49 26</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-49.5,-1511.5,-49.5,-1284.5</points>
<intersection>-1511.5 29</intersection>
<intersection>-1284.5 27</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>-49.5,-1511.5,184.5,-1511.5</points>
<connection>
<GID>659</GID>
<name>IN_1</name></connection>
<intersection>-49.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-440,8,-79</points>
<intersection>-440 14</intersection>
<intersection>-313.5 12</intersection>
<intersection>-153 5</intersection>
<intersection>-90.5 10</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-79,8,-79</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>8,-153,151,-153</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>8,-90.5,59.5,-90.5</points>
<connection>
<GID>390</GID>
<name>IN_4</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>8,-313.5,149.5,-313.5</points>
<connection>
<GID>532</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>8,-440,160.5,-440</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection>
<intersection>8.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>8.5,-622,8.5,-440</points>
<intersection>-622 16</intersection>
<intersection>-440 14</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>8.5,-622,168.5,-622</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>8.5 15</intersection>
<intersection>9 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>9,-1277,9,-622</points>
<intersection>-1277 22</intersection>
<intersection>-1043 20</intersection>
<intersection>-821 18</intersection>
<intersection>-622 16</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>9,-821,179,-821</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>9 17</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>9,-1043,172.5,-1043</points>
<connection>
<GID>576</GID>
<name>IN_1</name></connection>
<intersection>9 17</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>9,-1277,174.5,-1277</points>
<connection>
<GID>618</GID>
<name>IN_1</name></connection>
<intersection>9 17</intersection>
<intersection>9.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>9.5,-1504,9.5,-1277</points>
<intersection>-1504 24</intersection>
<intersection>-1277 22</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>9.5,-1504,183.5,-1504</points>
<connection>
<GID>660</GID>
<name>IN_1</name></connection>
<intersection>9.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>51,-305,51,-79.5</points>
<intersection>-305 18</intersection>
<intersection>-145.5 10</intersection>
<intersection>-89.5 16</intersection>
<intersection>-79.5 13</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>51,-145.5,150,-145.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>51 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>44,-79.5,51,-79.5</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<intersection>51 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>51,-89.5,59.5,-89.5</points>
<connection>
<GID>390</GID>
<name>IN_5</name></connection>
<intersection>51 3</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>51,-305,149.5,-305</points>
<connection>
<GID>533</GID>
<name>IN_1</name></connection>
<intersection>51 3</intersection>
<intersection>51.5 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>51.5,-1035.5,51.5,-305</points>
<intersection>-1035.5 26</intersection>
<intersection>-813.5 24</intersection>
<intersection>-614.5 22</intersection>
<intersection>-432.5 20</intersection>
<intersection>-305 18</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>51.5,-432.5,159.5,-432.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>51.5 19</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>51.5,-614.5,167.5,-614.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>51.5 19</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>51.5,-813.5,178,-813.5</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>51.5 19</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>51.5,-1035.5,171.5,-1035.5</points>
<connection>
<GID>577</GID>
<name>IN_1</name></connection>
<intersection>51.5 19</intersection>
<intersection>52 27</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>52,-1496.5,52,-1035.5</points>
<intersection>-1496.5 30</intersection>
<intersection>-1269.5 28</intersection>
<intersection>-1035.5 26</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>52,-1269.5,173.5,-1269.5</points>
<connection>
<GID>619</GID>
<name>IN_1</name></connection>
<intersection>52 27</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>52,-1496.5,182.5,-1496.5</points>
<connection>
<GID>661</GID>
<name>IN_1</name></connection>
<intersection>52 27</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-178,-35,-178,-22.5</points>
<intersection>-35 8</intersection>
<intersection>-22.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-186.5,-22.5,-178,-22.5</points>
<intersection>-186.5 9</intersection>
<intersection>-178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-178,-35,-175,-35</points>
<connection>
<GID>355</GID>
<name>J</name></connection>
<intersection>-178 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-186.5,-23,-186.5,-11</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-22.5 6</intersection>
<intersection>-11 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-227.5,-11,-186.5,-11</points>
<intersection>-227.5 14</intersection>
<intersection>-186.5 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-227.5,-14.5,-227.5,-11</points>
<intersection>-14.5 15</intersection>
<intersection>-11 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-238,-14.5,-227.5,-14.5</points>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<intersection>-227.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-193,-15.5,5,-15.5</points>
<intersection>-193 7</intersection>
<intersection>-137.5 6</intersection>
<intersection>-101 10</intersection>
<intersection>-72.5 12</intersection>
<intersection>-42.5 14</intersection>
<intersection>5 16</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-137.5,-20.5,-137.5,-15.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>-15.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-193,-22.5,-193,-15.5</points>
<intersection>-22.5 20</intersection>
<intersection>-15.5 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-101,-20,-101,-15.5</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>-15.5 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-72.5,-20.5,-72.5,-15.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>-15.5 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-42.5,-20.5,-42.5,-15.5</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>-15.5 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>5,-18.5,5,-15.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-223.5,-22.5,-188.5,-22.5</points>
<intersection>-223.5 23</intersection>
<intersection>-193 7</intersection>
<intersection>-188.5 26</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-223.5,-158,-223.5,-22.5</points>
<intersection>-158 24</intersection>
<intersection>-22.5 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-223.5,-158,-159.5,-158</points>
<intersection>-223.5 23</intersection>
<intersection>-159.5 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-159.5,-158,-159.5,-157</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>-158 24</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-188.5,-23,-188.5,-22.5</points>
<connection>
<GID>402</GID>
<name>IN_1</name></connection>
<intersection>-22.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-187.5,-39,-187.5,-29</points>
<connection>
<GID>402</GID>
<name>OUT</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-187.5,-39,-175,-39</points>
<connection>
<GID>355</GID>
<name>K</name></connection>
<intersection>-187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-139,-129,-139,-117.5</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>-117.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-144,-117.5,-144,-112</points>
<connection>
<GID>411</GID>
<name>OUT_0</name></connection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-144,-117.5,-139,-117.5</points>
<intersection>-144 1</intersection>
<intersection>-139 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-137,-129,-137,-117.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-117.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-131.5,-117.5,-131.5,-113</points>
<connection>
<GID>412</GID>
<name>OUT_0</name></connection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-137,-117.5,-131.5,-117.5</points>
<intersection>-137 0</intersection>
<intersection>-131.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-160.5,-151,-160.5,-138.5</points>
<connection>
<GID>409</GID>
<name>IN_2</name></connection>
<intersection>-138.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-138,-138.5,-138,-135</points>
<connection>
<GID>396</GID>
<name>OUT</name></connection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-160.5,-138.5,-138,-138.5</points>
<intersection>-160.5 0</intersection>
<intersection>-138 1</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-115.5,-63,-113.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>-113.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-60.5,-113.5,-60.5,-112</points>
<connection>
<GID>414</GID>
<name>OUT_0</name></connection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-63,-113.5,-60.5,-113.5</points>
<intersection>-63 0</intersection>
<intersection>-60.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-115.5,-65,-113.5</points>
<connection>
<GID>399</GID>
<name>IN_1</name></connection>
<intersection>-113.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-67.5,-113.5,-67.5,-112</points>
<connection>
<GID>413</GID>
<name>OUT_0</name></connection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-67.5,-113.5,-65,-113.5</points>
<intersection>-67.5 1</intersection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-158.5,-151,-158.5,-140.5</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>-140.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-64,-140.5,-64,-121.5</points>
<connection>
<GID>399</GID>
<name>OUT</name></connection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-158.5,-140.5,-64,-140.5</points>
<intersection>-158.5 0</intersection>
<intersection>-64 1</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.57746e-008,-114,-3.57746e-008,-112.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>-112.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>2.5,-112.5,2.5,-111</points>
<connection>
<GID>417</GID>
<name>OUT_0</name></connection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-3.57746e-008,-112.5,2.5,-112.5</points>
<intersection>-3.57746e-008 0</intersection>
<intersection>2.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-114,-2,-112.5</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<intersection>-112.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-3,-112.5,-3,-111.5</points>
<connection>
<GID>416</GID>
<name>OUT_0</name></connection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-3,-112.5,-2,-112.5</points>
<intersection>-3 1</intersection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-156.5,-151,-156.5,-143</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>-143 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1,-143,-1,-120</points>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<intersection>-143 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-156.5,-143,-1,-143</points>
<intersection>-156.5 0</intersection>
<intersection>-1 1</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-128,-37.5,-128,-20</points>
<intersection>-37.5 2</intersection>
<intersection>-35.5 1</intersection>
<intersection>-20 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-128,-35.5,-125.5,-35.5</points>
<connection>
<GID>357</GID>
<name>J</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-138.5,-37.5,-128,-37.5</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-135.5,-20,-128,-20</points>
<intersection>-135.5 4</intersection>
<intersection>-128 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-135.5,-20.5,-135.5,-20</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-20 3</intersection></vsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-136.5,-39.5,-136.5,-26.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-136.5,-39.5,-125.5,-39.5</points>
<connection>
<GID>357</GID>
<name>K</name></connection>
<intersection>-136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-35,-100,-26</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-100,-35,-99.5,-35</points>
<connection>
<GID>359</GID>
<name>J</name></connection>
<intersection>-100 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,-27.5,-92.5,-20</points>
<intersection>-27.5 1</intersection>
<intersection>-20 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-102,-27.5,-92.5,-27.5</points>
<intersection>-102 4</intersection>
<intersection>-92.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-99,-20,-92.5,-20</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>-92.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-102,-39,-102,-27.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>-39 6</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-102,-39,-99.5,-39</points>
<connection>
<GID>359</GID>
<name>K</name></connection>
<intersection>-102 4</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-73.5,-28,-67,-28</points>
<intersection>-73.5 3</intersection>
<intersection>-67 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-73.5,-37,-73.5,-28</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>-35.5 7</intersection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-67,-28,-67,-20.5</points>
<intersection>-28 1</intersection>
<intersection>-20.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-70.5,-20.5,-67,-20.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>-67 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-35.5,-69.5,-35.5</points>
<connection>
<GID>361</GID>
<name>J</name></connection>
<intersection>-73.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71.5,-39.5,-71.5,-26.5</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-39.5,-69.5,-39.5</points>
<connection>
<GID>361</GID>
<name>K</name></connection>
<intersection>-71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44.5,-37.5,-31,-37.5</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<connection>
<GID>363</GID>
<name>J</name></connection>
<intersection>-35 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-35,-37.5,-35,-19.5</points>
<intersection>-37.5 1</intersection>
<intersection>-19.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-40.5,-19.5,-35,-19.5</points>
<intersection>-40.5 6</intersection>
<intersection>-35 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-40.5,-20.5,-40.5,-19.5</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>-19.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-41.5,-41.5,-26.5</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41.5,-41.5,-31,-41.5</points>
<connection>
<GID>363</GID>
<name>K</name></connection>
<intersection>-41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-38,17.5,-38</points>
<connection>
<GID>385</GID>
<name>OUT</name></connection>
<connection>
<GID>365</GID>
<name>J</name></connection>
<intersection>10.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10.5,-38,10.5,-17</points>
<intersection>-38 1</intersection>
<intersection>-17 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>7,-17,10.5,-17</points>
<intersection>7 15</intersection>
<intersection>10.5 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>7,-18.5,7,-17</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>-17 8</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-42,6,-24.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-42,17.5,-42</points>
<connection>
<GID>365</GID>
<name>K</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-248,-8.5,-239,-8.5</points>
<connection>
<GID>420</GID>
<name>IN_1</name></connection>
<connection>
<GID>523</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-237,-8.5,-237,-7.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-231,-7.5,-231,-6</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-237,-7.5,-231,-7.5</points>
<intersection>-237 0</intersection>
<intersection>-231 1</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-252,-58,-252,-33</points>
<intersection>-58 1</intersection>
<intersection>-33 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-279.5,-58,-247.5,-58</points>
<connection>
<GID>393</GID>
<name>IN_1</name></connection>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<intersection>-252 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-252,-33,-246.5,-33</points>
<intersection>-252 0</intersection>
<intersection>-246.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-246.5,-41.5,-246.5,-33</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-33 4</intersection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-265.5,-56,-265.5,-40</points>
<intersection>-56 3</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-281,-40,-264,-40</points>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection>
<intersection>-265.5 0</intersection>
<intersection>-264 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-265.5,-56,-247.5,-56</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>-265.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-264,-40.5,-264,-40</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<intersection>-40 1</intersection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-248.5,-41.5,-248.5,-40.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-260,-40.5,-248.5,-40.5</points>
<connection>
<GID>395</GID>
<name>OUT_0</name></connection>
<intersection>-248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-247.5,-48,-242,-48</points>
<intersection>-247.5 5</intersection>
<intersection>-242 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-242,-48,-242,-43.5</points>
<intersection>-48 1</intersection>
<intersection>-43.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-247.5,-48,-247.5,-47.5</points>
<connection>
<GID>397</GID>
<name>OUT</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-242,-43.5,-238.5,-43.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-242 2</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-228,-43.5,-228,-27</points>
<intersection>-43.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-232.5,-43.5,-228,-43.5</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<intersection>-228 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-228,-27,-158.5,-27</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>-228 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-232.5,-46.5,-159.5,-46.5</points>
<connection>
<GID>388</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>-205 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-205,-151,-205,-46.5</points>
<intersection>-151 8</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-205,-151,-162.5,-151</points>
<connection>
<GID>409</GID>
<name>IN_3</name></connection>
<intersection>-205 7</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-241.5,138.5,401.5,138.5</points>
<intersection>-241.5 15</intersection>
<intersection>-234 16</intersection>
<intersection>401.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>401.5,-250,401.5,138.5</points>
<intersection>-250 3</intersection>
<intersection>138.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>244.5,-250,401.5,-250</points>
<intersection>244.5 14</intersection>
<intersection>260.5 13</intersection>
<intersection>274 12</intersection>
<intersection>289 11</intersection>
<intersection>299.5 10</intersection>
<intersection>312.5 9</intersection>
<intersection>401.5 2</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>312.5,-250,312.5,-238.5</points>
<connection>
<GID>422</GID>
<name>clock</name></connection>
<intersection>-250 3</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>299.5,-250,299.5,-238.5</points>
<connection>
<GID>415</GID>
<name>clock</name></connection>
<intersection>-250 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>289,-250,289,-238.5</points>
<connection>
<GID>410</GID>
<name>clock</name></connection>
<intersection>-250 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>274,-250,274,-238.5</points>
<connection>
<GID>403</GID>
<name>clock</name></connection>
<intersection>-250 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>260.5,-250,260.5,-238.5</points>
<connection>
<GID>394</GID>
<name>clock</name></connection>
<intersection>-250 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>244.5,-293,244.5,-238</points>
<connection>
<GID>368</GID>
<name>clock</name></connection>
<intersection>-293 196</intersection>
<intersection>-250 3</intersection>
<intersection>-238 17</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-241.5,138.5,-241.5,149</points>
<connection>
<GID>473</GID>
<name>CLK</name></connection>
<intersection>138.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-234,138.5,-234,149</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>138.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>109,-238,244.5,-238</points>
<intersection>109 18</intersection>
<intersection>215 210</intersection>
<intersection>244.5 14</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>109,-363,109,-238</points>
<intersection>-363 41</intersection>
<intersection>-238 17</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>108.5,-363,311,-363</points>
<connection>
<GID>334</GID>
<name>clock</name></connection>
<intersection>108.5 89</intersection>
<intersection>109 18</intersection>
<intersection>213.5 215</intersection>
<intersection>244 52</intersection>
<intersection>259.5 51</intersection>
<intersection>273 50</intersection>
<intersection>287 49</intersection>
<intersection>298 48</intersection>
<intersection>311 47</intersection></hsegment>
<vsegment>
<ID>47</ID>
<points>311,-363.5,311,-363</points>
<intersection>-363.5 88</intersection>
<intersection>-363 41</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>298,-363.5,298,-363</points>
<intersection>-363.5 87</intersection>
<intersection>-363 41</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>287,-363.5,287,-363</points>
<intersection>-363.5 86</intersection>
<intersection>-363 41</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>273,-363.5,273,-363</points>
<intersection>-363.5 85</intersection>
<intersection>-363 41</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>259.5,-363.5,259.5,-363</points>
<intersection>-363.5 84</intersection>
<intersection>-363 41</intersection></vsegment>
<vsegment>
<ID>52</ID>
<points>244,-410,244,-363</points>
<intersection>-410 198</intersection>
<intersection>-363 41</intersection></vsegment>
<hsegment>
<ID>84</ID>
<points>259.5,-363.5,260,-363.5</points>
<connection>
<GID>75</GID>
<name>clock</name></connection>
<intersection>259.5 51</intersection></hsegment>
<hsegment>
<ID>85</ID>
<points>273,-363.5,273.5,-363.5</points>
<connection>
<GID>88</GID>
<name>clock</name></connection>
<intersection>273 50</intersection></hsegment>
<hsegment>
<ID>86</ID>
<points>287,-363.5,288.5,-363.5</points>
<connection>
<GID>92</GID>
<name>clock</name></connection>
<intersection>287 49</intersection></hsegment>
<hsegment>
<ID>87</ID>
<points>298,-363.5,299,-363.5</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>298 48</intersection></hsegment>
<hsegment>
<ID>88</ID>
<points>311,-363.5,312,-363.5</points>
<connection>
<GID>98</GID>
<name>clock</name></connection>
<intersection>311 47</intersection></hsegment>
<vsegment>
<ID>89</ID>
<points>108.5,-918,108.5,-363</points>
<intersection>-918 109</intersection>
<intersection>-916.5 138</intersection>
<intersection>-706.5 122</intersection>
<intersection>-537 93</intersection>
<intersection>-363 41</intersection></vsegment>
<hsegment>
<ID>93</ID>
<points>108.5,-537,322,-537</points>
<intersection>108.5 89</intersection>
<intersection>189.5 213</intersection>
<intersection>254 104</intersection>
<intersection>270 103</intersection>
<intersection>283.5 102</intersection>
<intersection>298.5 101</intersection>
<intersection>309 100</intersection>
<intersection>322 99</intersection></hsegment>
<vsegment>
<ID>99</ID>
<points>322,-537,322,-525.5</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>-537 93</intersection></vsegment>
<vsegment>
<ID>100</ID>
<points>309,-537,309,-525.5</points>
<connection>
<GID>31</GID>
<name>clock</name></connection>
<intersection>-537 93</intersection></vsegment>
<vsegment>
<ID>101</ID>
<points>298.5,-537,298.5,-525.5</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>-537 93</intersection></vsegment>
<vsegment>
<ID>102</ID>
<points>283.5,-537,283.5,-525.5</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-537 93</intersection></vsegment>
<vsegment>
<ID>103</ID>
<points>270,-537,270,-525.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>-537 93</intersection></vsegment>
<vsegment>
<ID>104</ID>
<points>254,-579,254,-525</points>
<connection>
<GID>147</GID>
<name>clock</name></connection>
<intersection>-579 200</intersection>
<intersection>-537 93</intersection></vsegment>
<hsegment>
<ID>109</ID>
<points>108,-918,340.5,-918</points>
<intersection>108 153</intersection>
<intersection>108.5 89</intersection>
<intersection>204.5 219</intersection>
<intersection>272.5 205</intersection>
<intersection>288.5 119</intersection>
<intersection>302 118</intersection>
<intersection>317 117</intersection>
<intersection>327.5 116</intersection>
<intersection>340.5 115</intersection></hsegment>
<vsegment>
<ID>115</ID>
<points>340.5,-918,340.5,-906.5</points>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<intersection>-918 109</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>327.5,-918,327.5,-906.5</points>
<connection>
<GID>282</GID>
<name>clock</name></connection>
<intersection>-918 109</intersection></vsegment>
<vsegment>
<ID>117</ID>
<points>317,-918,317,-906.5</points>
<connection>
<GID>281</GID>
<name>clock</name></connection>
<intersection>-918 109</intersection></vsegment>
<vsegment>
<ID>118</ID>
<points>302,-918,302,-906.5</points>
<connection>
<GID>280</GID>
<name>clock</name></connection>
<intersection>-918 109</intersection></vsegment>
<vsegment>
<ID>119</ID>
<points>288.5,-918,288.5,-906.5</points>
<connection>
<GID>279</GID>
<name>clock</name></connection>
<intersection>-918 109</intersection></vsegment>
<hsegment>
<ID>122</ID>
<points>108.5,-706.5,262,-706.5</points>
<intersection>108.5 89</intersection>
<intersection>191 221</intersection>
<intersection>262 137</intersection></hsegment>
<hsegment>
<ID>126</ID>
<points>262,-719,330,-719</points>
<intersection>262 137</intersection>
<intersection>278 136</intersection>
<intersection>291.5 135</intersection>
<intersection>306.5 134</intersection>
<intersection>317 133</intersection>
<intersection>330 132</intersection></hsegment>
<vsegment>
<ID>132</ID>
<points>330,-719,330,-707.5</points>
<connection>
<GID>200</GID>
<name>clock</name></connection>
<intersection>-719 126</intersection></vsegment>
<vsegment>
<ID>133</ID>
<points>317,-719,317,-707.5</points>
<connection>
<GID>199</GID>
<name>clock</name></connection>
<intersection>-719 126</intersection></vsegment>
<vsegment>
<ID>134</ID>
<points>306.5,-719,306.5,-707.5</points>
<connection>
<GID>198</GID>
<name>clock</name></connection>
<intersection>-719 126</intersection></vsegment>
<vsegment>
<ID>135</ID>
<points>291.5,-719,291.5,-707.5</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>-719 126</intersection></vsegment>
<vsegment>
<ID>136</ID>
<points>278,-719,278,-707.5</points>
<connection>
<GID>196</GID>
<name>clock</name></connection>
<intersection>-719 126</intersection></vsegment>
<vsegment>
<ID>137</ID>
<points>262,-764.5,262,-706.5</points>
<connection>
<GID>278</GID>
<name>clock</name></connection>
<intersection>-764.5 227</intersection>
<intersection>-719 126</intersection>
<intersection>-706.5 122</intersection></vsegment>
<hsegment>
<ID>138</ID>
<points>108,-916.5,108.5,-916.5</points>
<intersection>108 153</intersection>
<intersection>108.5 89</intersection></hsegment>
<hsegment>
<ID>142</ID>
<points>108,-1140,334,-1140</points>
<intersection>108 153</intersection>
<intersection>207.5 218</intersection>
<intersection>266 194</intersection>
<intersection>282 152</intersection>
<intersection>295.5 151</intersection>
<intersection>310.5 150</intersection>
<intersection>321 149</intersection>
<intersection>334 148</intersection></hsegment>
<vsegment>
<ID>148</ID>
<points>334,-1140,334,-1128.5</points>
<connection>
<GID>335</GID>
<name>clock</name></connection>
<intersection>-1140 142</intersection></vsegment>
<vsegment>
<ID>149</ID>
<points>321,-1140,321,-1128.5</points>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<intersection>-1140 142</intersection></vsegment>
<vsegment>
<ID>150</ID>
<points>310.5,-1140,310.5,-1128.5</points>
<connection>
<GID>323</GID>
<name>clock</name></connection>
<intersection>-1140 142</intersection></vsegment>
<vsegment>
<ID>151</ID>
<points>295.5,-1140,295.5,-1128.5</points>
<intersection>-1140 142</intersection>
<intersection>-1128.5 217</intersection></vsegment>
<vsegment>
<ID>152</ID>
<points>282,-1140,282,-1128.5</points>
<connection>
<GID>321</GID>
<name>clock</name></connection>
<intersection>-1140 142</intersection></vsegment>
<vsegment>
<ID>153</ID>
<points>108,-1601,108,-916.5</points>
<intersection>-1601 174</intersection>
<intersection>-1589 192</intersection>
<intersection>-1420.5 208</intersection>
<intersection>-1374 158</intersection>
<intersection>-1140 142</intersection>
<intersection>-961 204</intersection>
<intersection>-918 109</intersection>
<intersection>-916.5 138</intersection></vsegment>
<hsegment>
<ID>158</ID>
<points>108,-1374,336,-1374</points>
<intersection>108 153</intersection>
<intersection>207.5 222</intersection>
<intersection>268 169</intersection>
<intersection>284 168</intersection>
<intersection>297.5 167</intersection>
<intersection>312.5 166</intersection>
<intersection>323 209</intersection>
<intersection>336 164</intersection></hsegment>
<vsegment>
<ID>164</ID>
<points>336,-1374,336,-1362.5</points>
<connection>
<GID>583</GID>
<name>clock</name></connection>
<intersection>-1374 158</intersection></vsegment>
<vsegment>
<ID>166</ID>
<points>312.5,-1374,312.5,-1362.5</points>
<connection>
<GID>581</GID>
<name>clock</name></connection>
<intersection>-1374 158</intersection></vsegment>
<vsegment>
<ID>167</ID>
<points>297.5,-1374,297.5,-1362.5</points>
<connection>
<GID>580</GID>
<name>clock</name></connection>
<intersection>-1374 158</intersection></vsegment>
<vsegment>
<ID>168</ID>
<points>284,-1374,284,-1362.5</points>
<connection>
<GID>579</GID>
<name>clock</name></connection>
<intersection>-1374 158</intersection></vsegment>
<vsegment>
<ID>169</ID>
<points>268,-1374,268,-1362</points>
<connection>
<GID>620</GID>
<name>clock</name></connection>
<intersection>-1374 158</intersection></vsegment>
<hsegment>
<ID>174</ID>
<points>108,-1601,345,-1601</points>
<intersection>108 153</intersection>
<intersection>228.5 224</intersection>
<intersection>293 184</intersection>
<intersection>306.5 183</intersection>
<intersection>321.5 182</intersection>
<intersection>332 181</intersection>
<intersection>345 180</intersection></hsegment>
<vsegment>
<ID>180</ID>
<points>345,-1601,345,-1589.5</points>
<connection>
<GID>625</GID>
<name>clock</name></connection>
<intersection>-1601 174</intersection></vsegment>
<vsegment>
<ID>181</ID>
<points>332,-1601,332,-1589.5</points>
<connection>
<GID>624</GID>
<name>clock</name></connection>
<intersection>-1601 174</intersection></vsegment>
<vsegment>
<ID>182</ID>
<points>321.5,-1601,321.5,-1589.5</points>
<connection>
<GID>623</GID>
<name>clock</name></connection>
<intersection>-1601 174</intersection></vsegment>
<vsegment>
<ID>183</ID>
<points>306.5,-1601,306.5,-1589.5</points>
<connection>
<GID>622</GID>
<name>clock</name></connection>
<intersection>-1601 174</intersection></vsegment>
<vsegment>
<ID>184</ID>
<points>293,-1601,293,-1589.5</points>
<connection>
<GID>621</GID>
<name>clock</name></connection>
<intersection>-1601 174</intersection></vsegment>
<hsegment>
<ID>192</ID>
<points>108,-1589,277,-1589</points>
<connection>
<GID>662</GID>
<name>clock</name></connection>
<intersection>108 153</intersection></hsegment>
<vsegment>
<ID>194</ID>
<points>266,-1186,266,-1128</points>
<connection>
<GID>578</GID>
<name>clock</name></connection>
<intersection>-1186 229</intersection>
<intersection>-1140 142</intersection></vsegment>
<hsegment>
<ID>196</ID>
<points>244.5,-293,311.5,-293</points>
<connection>
<GID>2090</GID>
<name>clock</name></connection>
<intersection>244.5 14</intersection></hsegment>
<hsegment>
<ID>198</ID>
<points>244,-410,302,-410</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>244 52</intersection></hsegment>
<hsegment>
<ID>200</ID>
<points>254,-579,308,-579</points>
<connection>
<GID>55</GID>
<name>clock</name></connection>
<intersection>254 104</intersection></hsegment>
<hsegment>
<ID>204</ID>
<points>108,-961,324,-961</points>
<connection>
<GID>188</GID>
<name>clock</name></connection>
<intersection>108 153</intersection></hsegment>
<vsegment>
<ID>205</ID>
<points>272.5,-918,272.5,-906</points>
<connection>
<GID>320</GID>
<name>clock</name></connection>
<intersection>-918 109</intersection></vsegment>
<hsegment>
<ID>208</ID>
<points>108,-1420.5,323,-1420.5</points>
<connection>
<GID>267</GID>
<name>clock</name></connection>
<intersection>108 153</intersection></hsegment>
<vsegment>
<ID>209</ID>
<points>323,-1374,323,-1362.5</points>
<connection>
<GID>582</GID>
<name>clock</name></connection>
<intersection>-1374 158</intersection></vsegment>
<vsegment>
<ID>210</ID>
<points>215,-254.5,215,-238</points>
<intersection>-254.5 211</intersection>
<intersection>-238 17</intersection></vsegment>
<hsegment>
<ID>211</ID>
<points>215,-254.5,219,-254.5</points>
<connection>
<GID>1783</GID>
<name>clock</name></connection>
<intersection>215 210</intersection></hsegment>
<vsegment>
<ID>213</ID>
<points>189.5,-550,189.5,-537</points>
<intersection>-550 214</intersection>
<intersection>-537 93</intersection></vsegment>
<hsegment>
<ID>214</ID>
<points>189.5,-550,192,-550</points>
<connection>
<GID>1808</GID>
<name>clock</name></connection>
<intersection>189.5 213</intersection></hsegment>
<vsegment>
<ID>215</ID>
<points>213.5,-379,213.5,-363</points>
<intersection>-379 216</intersection>
<intersection>-363 41</intersection></vsegment>
<hsegment>
<ID>216</ID>
<points>213.5,-379,216,-379</points>
<connection>
<GID>1796</GID>
<name>clock</name></connection>
<intersection>213.5 215</intersection></hsegment>
<hsegment>
<ID>217</ID>
<points>295.5,-1128.5,296,-1128.5</points>
<connection>
<GID>322</GID>
<name>clock</name></connection>
<intersection>295.5 151</intersection></hsegment>
<vsegment>
<ID>218</ID>
<points>207.5,-1149,207.5,-1140</points>
<connection>
<GID>54</GID>
<name>clock</name></connection>
<intersection>-1140 142</intersection></vsegment>
<vsegment>
<ID>219</ID>
<points>204.5,-926,204.5,-918</points>
<intersection>-926 220</intersection>
<intersection>-918 109</intersection></vsegment>
<hsegment>
<ID>220</ID>
<points>204.5,-926,209,-926</points>
<connection>
<GID>40</GID>
<name>clock</name></connection>
<intersection>204.5 219</intersection></hsegment>
<vsegment>
<ID>221</ID>
<points>191,-717.5,191,-706.5</points>
<connection>
<GID>15</GID>
<name>clock</name></connection>
<intersection>-706.5 122</intersection></vsegment>
<vsegment>
<ID>222</ID>
<points>207.5,-1382.5,207.5,-1374</points>
<intersection>-1382.5 223</intersection>
<intersection>-1374 158</intersection></vsegment>
<hsegment>
<ID>223</ID>
<points>207.5,-1382.5,209.5,-1382.5</points>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<intersection>207.5 222</intersection></hsegment>
<vsegment>
<ID>224</ID>
<points>228.5,-1611,228.5,-1601</points>
<intersection>-1611 225</intersection>
<intersection>-1601 174</intersection></vsegment>
<hsegment>
<ID>225</ID>
<points>228.5,-1611,232,-1611</points>
<connection>
<GID>177</GID>
<name>clock</name></connection>
<intersection>228.5 224</intersection></hsegment>
<hsegment>
<ID>227</ID>
<points>262,-764.5,316,-764.5</points>
<connection>
<GID>162</GID>
<name>clock</name></connection>
<intersection>262 137</intersection></hsegment>
<hsegment>
<ID>229</ID>
<points>266,-1186,318.5,-1186</points>
<connection>
<GID>242</GID>
<name>clock</name></connection>
<intersection>266 194</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,85.5,14,86.5</points>
<intersection>85.5 2</intersection>
<intersection>86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,86.5,14,86.5</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,85.5,19,85.5</points>
<connection>
<GID>431</GID>
<name>Q</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-217,98,-217,102.5</points>
<intersection>98 1</intersection>
<intersection>102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-220.5,98,-217,98</points>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>-217 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-217,102.5,-213.5,102.5</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>-217 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,-1133,330.5,-1125.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327,-1125.5,330.5,-1125.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-226.5,85.5,3.5,85.5</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<connection>
<GID>472</GID>
<name>clear</name></connection>
<connection>
<GID>466</GID>
<name>clear</name></connection>
<connection>
<GID>464</GID>
<name>clear</name></connection>
<connection>
<GID>462</GID>
<name>clear</name></connection>
<connection>
<GID>474</GID>
<name>clear</name></connection>
<intersection>-226.5 6</intersection>
<intersection>-90 4</intersection>
<intersection>-44.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-44.5,85,-44.5,85.5</points>
<connection>
<GID>469</GID>
<name>clear</name></connection>
<intersection>85.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-90,49.5,-90,85.5</points>
<intersection>49.5 5</intersection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-90,49.5,1,49.5</points>
<intersection>-90 4</intersection>
<intersection>-81 13</intersection>
<intersection>-64.5 12</intersection>
<intersection>-50 11</intersection>
<intersection>-33 10</intersection>
<intersection>-17 9</intersection>
<intersection>1 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-226.5,85.5,-226.5,105.5</points>
<intersection>85.5 1</intersection>
<intersection>105.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-227,105.5,-226.5,105.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>-226.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>1,49.5,1,50.5</points>
<connection>
<GID>492</GID>
<name>clear</name></connection>
<intersection>49.5 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-17,49.5,-17,50.5</points>
<connection>
<GID>491</GID>
<name>clear</name></connection>
<intersection>49.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-33,49.5,-33,50.5</points>
<connection>
<GID>490</GID>
<name>clear</name></connection>
<intersection>49.5 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-50,49.5,-50,50.5</points>
<connection>
<GID>488</GID>
<name>clear</name></connection>
<intersection>49.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-64.5,49.5,-64.5,50.5</points>
<connection>
<GID>487</GID>
<name>clear</name></connection>
<intersection>49.5 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-81,49.5,-81,50.5</points>
<connection>
<GID>485</GID>
<name>clear</name></connection>
<intersection>49.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-220.5,96,-180.5,96</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>-180.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-180.5,94,-180.5,96</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<intersection>96 1</intersection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-239,106.5,-239,110.5</points>
<intersection>106.5 2</intersection>
<intersection>110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-245.5,110.5,-239,110.5</points>
<connection>
<GID>454</GID>
<name>IN_1</name></connection>
<intersection>-239 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-239,106.5,-233,106.5</points>
<connection>
<GID>452</GID>
<name>OUT</name></connection>
<intersection>-239 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,89.5,7,172.5</points>
<intersection>89.5 2</intersection>
<intersection>172.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-89.5,172.5,7,172.5</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,89.5,19,89.5</points>
<connection>
<GID>431</GID>
<name>nQ</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-218.5,158.5,-173,158.5</points>
<connection>
<GID>453</GID>
<name>clear</name></connection>
<connection>
<GID>451</GID>
<name>clear</name></connection>
<connection>
<GID>450</GID>
<name>clear</name></connection>
<intersection>-218.5 13</intersection>
<intersection>-173 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-173,157.5,-173,158.5</points>
<connection>
<GID>455</GID>
<name>clear</name></connection>
<intersection>157.5 5</intersection>
<intersection>158.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-173,157.5,-91.5,157.5</points>
<connection>
<GID>458</GID>
<name>clear</name></connection>
<connection>
<GID>457</GID>
<name>clear</name></connection>
<intersection>-173 4</intersection>
<intersection>-110.5 12</intersection>
<intersection>-91.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-91.5,150.5,-91.5,157.5</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>157.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-110.5,157.5,-110.5,164.5</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<intersection>157.5 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-218.5,123.5,-218.5,158.5</points>
<intersection>123.5 14</intersection>
<intersection>158.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-218.5,123.5,-127.5,123.5</points>
<connection>
<GID>507</GID>
<name>clear</name></connection>
<connection>
<GID>505</GID>
<name>clear</name></connection>
<connection>
<GID>503</GID>
<name>clear</name></connection>
<connection>
<GID>500</GID>
<name>clear</name></connection>
<connection>
<GID>499</GID>
<name>clear</name></connection>
<connection>
<GID>495</GID>
<name>clear</name></connection>
<intersection>-218.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122.5,177,-89.5,177</points>
<intersection>-122.5 3</intersection>
<intersection>-89.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122.5,173,-122.5,177</points>
<intersection>173 5</intersection>
<intersection>177 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-89.5,174.5,-89.5,177</points>
<connection>
<GID>438</GID>
<name>IN_1</name></connection>
<intersection>177 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-123.5,173,-122.5,173</points>
<connection>
<GID>489</GID>
<name>OUT</name></connection>
<intersection>-122.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343.5,-1132.5,343.5,-1125.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>-1125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>340,-1125.5,343.5,-1125.5</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>343.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-1142.5,276,-1137</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>-1142.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>291,-1148.5,291,-1142.5</points>
<connection>
<GID>419</GID>
<name>IN_3</name></connection>
<intersection>-1142.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>276,-1142.5,291,-1142.5</points>
<intersection>276 0</intersection>
<intersection>291 1</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-238,97,-226.5,97</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<connection>
<GID>449</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-244,98,-244,108.5</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-245.5,108.5,-244,108.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-244 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-259.5,109.5,-251.5,109.5</points>
<connection>
<GID>468</GID>
<name>N_in1</name></connection>
<connection>
<GID>454</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,165.5,-100,173.5</points>
<intersection>165.5 1</intersection>
<intersection>173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-104.5,165.5,-100,165.5</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-100,173.5,-95.5,173.5</points>
<connection>
<GID>438</GID>
<name>OUT</name></connection>
<intersection>-100 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,79.5,-100,163.5</points>
<intersection>79.5 3</intersection>
<intersection>163.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-104.5,163.5,-100,163.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>-100 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-242,79.5,9.5,79.5</points>
<connection>
<GID>447</GID>
<name>OUT_0</name></connection>
<intersection>-100 0</intersection>
<intersection>9.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>9.5,79.5,9.5,84.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>79.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-193.5,160.5,-193.5,173</points>
<intersection>160.5 4</intersection>
<intersection>164.5 2</intersection>
<intersection>173 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-195,173,-184,173</points>
<connection>
<GID>476</GID>
<name>OUT</name></connection>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>-193.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-193.5,164.5,-192,164.5</points>
<connection>
<GID>453</GID>
<name>J</name></connection>
<intersection>-193.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-193.5,160.5,-192,160.5</points>
<connection>
<GID>453</GID>
<name>K</name></connection>
<intersection>-193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-177,160,-177,172</points>
<intersection>160 4</intersection>
<intersection>164 2</intersection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-178,172,-169,172</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>-177 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-177,164,-176,164</points>
<connection>
<GID>455</GID>
<name>J</name></connection>
<intersection>-177 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-177,160,-176,160</points>
<connection>
<GID>455</GID>
<name>K</name></connection>
<intersection>-177 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-161.5,159.5,-161.5,171</points>
<intersection>159.5 4</intersection>
<intersection>163.5 2</intersection>
<intersection>171 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-163,171,-151.5,171</points>
<connection>
<GID>483</GID>
<name>OUT</name></connection>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-161.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-161.5,163.5,-160,163.5</points>
<connection>
<GID>457</GID>
<name>J</name></connection>
<intersection>-161.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-161.5,159.5,-160,159.5</points>
<connection>
<GID>457</GID>
<name>K</name></connection>
<intersection>-161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-144.5,159.5,-144.5,170</points>
<intersection>159.5 4</intersection>
<intersection>163.5 2</intersection>
<intersection>170 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-145.5,170,-144.5,170</points>
<connection>
<GID>486</GID>
<name>OUT</name></connection>
<intersection>-144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-144.5,163.5,-143,163.5</points>
<connection>
<GID>458</GID>
<name>J</name></connection>
<intersection>-144.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-144.5,159.5,-143,159.5</points>
<connection>
<GID>458</GID>
<name>K</name></connection>
<intersection>-144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-215.5,164.5,-208,164.5</points>
<connection>
<GID>450</GID>
<name>Q</name></connection>
<connection>
<GID>451</GID>
<name>J</name></connection>
<intersection>-214.5 3</intersection>
<intersection>-212 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-214.5,129.5,-214.5,164.5</points>
<intersection>129.5 10</intersection>
<intersection>145 4</intersection>
<intersection>160.5 9</intersection>
<intersection>164.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-214.5,145,-127.5,145</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-214.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-212,164.5,-212,174</points>
<intersection>164.5 1</intersection>
<intersection>174 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-212,174,-201,174</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>-212 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-214.5,160.5,-208,160.5</points>
<connection>
<GID>451</GID>
<name>K</name></connection>
<intersection>-214.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-214.5,129.5,-212.5,129.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>-214.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-227.5,155,38,155</points>
<intersection>-227.5 3</intersection>
<intersection>-212 4</intersection>
<intersection>-196 32</intersection>
<intersection>-195 5</intersection>
<intersection>-181.5 31</intersection>
<intersection>-179 16</intersection>
<intersection>-164.5 30</intersection>
<intersection>-162.5 15</intersection>
<intersection>-148.5 29</intersection>
<intersection>-147.5 18</intersection>
<intersection>-130.5 28</intersection>
<intersection>38 35</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-227.5,126.5,-227.5,162.5</points>
<intersection>126.5 33</intersection>
<intersection>150 39</intersection>
<intersection>155 1</intersection>
<intersection>162.5 13</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-212,155,-212,162.5</points>
<intersection>155 1</intersection>
<intersection>162.5 14</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-195,155,-195,162.5</points>
<intersection>155 1</intersection>
<intersection>162.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-195,162.5,-192,162.5</points>
<connection>
<GID>453</GID>
<name>clock</name></connection>
<intersection>-195 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-227.5,162.5,-221.5,162.5</points>
<connection>
<GID>450</GID>
<name>clock</name></connection>
<intersection>-227.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-212,162.5,-208,162.5</points>
<connection>
<GID>451</GID>
<name>clock</name></connection>
<intersection>-212 4</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-162.5,155,-162.5,161.5</points>
<intersection>155 1</intersection>
<intersection>161.5 21</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-179,155,-179,162</points>
<intersection>155 1</intersection>
<intersection>162 19</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-147.5,155,-147.5,161.5</points>
<intersection>155 1</intersection>
<intersection>161.5 20</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-179,162,-176,162</points>
<connection>
<GID>455</GID>
<name>clock</name></connection>
<intersection>-179 16</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-147.5,161.5,-143,161.5</points>
<connection>
<GID>458</GID>
<name>clock</name></connection>
<intersection>-147.5 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-162.5,161.5,-160,161.5</points>
<connection>
<GID>457</GID>
<name>clock</name></connection>
<intersection>-162.5 15</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-130.5,126.5,-130.5,155</points>
<connection>
<GID>507</GID>
<name>clock</name></connection>
<intersection>155 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>-148.5,126.5,-148.5,155</points>
<connection>
<GID>505</GID>
<name>clock</name></connection>
<intersection>155 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-164.5,126.5,-164.5,155</points>
<connection>
<GID>503</GID>
<name>clock</name></connection>
<intersection>155 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-181.5,126.5,-181.5,155</points>
<connection>
<GID>500</GID>
<name>clock</name></connection>
<intersection>155 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-196,126.5,-196,155</points>
<connection>
<GID>499</GID>
<name>clock</name></connection>
<intersection>155 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-227.5,126.5,-212.5,126.5</points>
<connection>
<GID>495</GID>
<name>clock</name></connection>
<intersection>-227.5 3</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>38,87.5,38,155</points>
<intersection>87.5 36</intersection>
<intersection>155 1</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>25,87.5,38,87.5</points>
<connection>
<GID>431</GID>
<name>clock</name></connection>
<intersection>38 35</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-228,150,-227.5,150</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<intersection>-227.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-201,129.5,-201,172</points>
<connection>
<GID>476</GID>
<name>IN_1</name></connection>
<intersection>129.5 8</intersection>
<intersection>146 1</intersection>
<intersection>164.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-201,146,-127.5,146</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>-201 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-202,164.5,-201,164.5</points>
<connection>
<GID>451</GID>
<name>Q</name></connection>
<intersection>-201 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-201,129.5,-196,129.5</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>-201 0</intersection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-169,148,-127.5,148</points>
<connection>
<GID>465</GID>
<name>IN_3</name></connection>
<intersection>-169 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-169,129.5,-169,174</points>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<intersection>129.5 9</intersection>
<intersection>148 1</intersection>
<intersection>164 4</intersection>
<intersection>174 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-170,164,-169,164</points>
<connection>
<GID>455</GID>
<name>Q</name></connection>
<intersection>-169 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-169,174,-129.5,174</points>
<connection>
<GID>489</GID>
<name>IN_1</name></connection>
<intersection>-169 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-169,129.5,-164.5,129.5</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>-169 3</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-185,129.5,-185,176</points>
<intersection>129.5 9</intersection>
<intersection>147 4</intersection>
<intersection>164.5 3</intersection>
<intersection>171 2</intersection>
<intersection>176 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-185,171,-184,171</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>-185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-186,164.5,-185,164.5</points>
<connection>
<GID>453</GID>
<name>Q</name></connection>
<intersection>-185 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-185,147,-127.5,147</points>
<connection>
<GID>465</GID>
<name>IN_2</name></connection>
<intersection>-185 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-185,176,-129.5,176</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>-185 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-185,129.5,-181.5,129.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-185 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-153,129.5,-153,172</points>
<intersection>129.5 8</intersection>
<intersection>149 3</intersection>
<intersection>163.5 1</intersection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-154,163.5,-153,163.5</points>
<connection>
<GID>457</GID>
<name>Q</name></connection>
<intersection>-153 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-153,172,-129.5,172</points>
<connection>
<GID>489</GID>
<name>IN_2</name></connection>
<intersection>-153 0</intersection>
<intersection>-151.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-153,149,-127.5,149</points>
<connection>
<GID>465</GID>
<name>IN_4</name></connection>
<intersection>-153 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-151.5,169,-151.5,172</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-153,129.5,-148.5,129.5</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>-153 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-135,129.5,-135,170</points>
<intersection>129.5 5</intersection>
<intersection>150 2</intersection>
<intersection>163.5 1</intersection>
<intersection>170 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-137,163.5,-135,163.5</points>
<connection>
<GID>458</GID>
<name>Q</name></connection>
<intersection>-135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-135,150,-127.5,150</points>
<connection>
<GID>465</GID>
<name>IN_5</name></connection>
<intersection>-135 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-135,170,-129.5,170</points>
<connection>
<GID>489</GID>
<name>IN_3</name></connection>
<intersection>-135 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-135,129.5,-130.5,129.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>-135 0</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-205,115,-112.5,115</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>-205 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-205,105.5,-205,129.5</points>
<intersection>105.5 8</intersection>
<intersection>115 1</intersection>
<intersection>129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-206.5,129.5,-205,129.5</points>
<connection>
<GID>495</GID>
<name>OUT_0</name></connection>
<intersection>-205 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-206.5,105.5,-205,105.5</points>
<connection>
<GID>448</GID>
<name>IN_3</name></connection>
<intersection>-205 3</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-188.5,116,-112.5,116</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<intersection>-188.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-188.5,103.5,-188.5,129.5</points>
<intersection>103.5 8</intersection>
<intersection>116 1</intersection>
<intersection>129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-190,129.5,-188.5,129.5</points>
<connection>
<GID>499</GID>
<name>OUT_0</name></connection>
<intersection>-188.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-206.5,103.5,-188.5,103.5</points>
<connection>
<GID>448</GID>
<name>IN_2</name></connection>
<intersection>-188.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-174.5,117,-112.5,117</points>
<connection>
<GID>509</GID>
<name>IN_2</name></connection>
<intersection>-174.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-174.5,101.5,-174.5,129.5</points>
<intersection>101.5 8</intersection>
<intersection>117 1</intersection>
<intersection>129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-175.5,129.5,-174.5,129.5</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<intersection>-174.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-206.5,101.5,-174.5,101.5</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>-174.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-156,118,-112.5,118</points>
<connection>
<GID>509</GID>
<name>IN_3</name></connection>
<intersection>-156 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-156,99.5,-156,129.5</points>
<intersection>99.5 8</intersection>
<intersection>118 1</intersection>
<intersection>129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-158.5,129.5,-156,129.5</points>
<connection>
<GID>503</GID>
<name>OUT_0</name></connection>
<intersection>-156 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-206.5,99.5,-156,99.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>-156 3</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-174.5,119,-112.5,119</points>
<connection>
<GID>509</GID>
<name>IN_4</name></connection>
<intersection>-174.5 7</intersection>
<intersection>-141.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-141.5,119,-141.5,129.5</points>
<intersection>119 1</intersection>
<intersection>129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-142.5,129.5,-141.5,129.5</points>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection>
<intersection>-141.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-174.5,95,-174.5,119</points>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>119 1</intersection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121.5,120,-112.5,120</points>
<connection>
<GID>509</GID>
<name>IN_5</name></connection>
<intersection>-121.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-121.5,93,-121.5,129.5</points>
<intersection>93 8</intersection>
<intersection>120 1</intersection>
<intersection>129.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-124.5,129.5,-121.5,129.5</points>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection>
<intersection>-121.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-174.5,93,-121.5,93</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>-121.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,87.5,-65,100</points>
<intersection>87.5 4</intersection>
<intersection>91.5 2</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,100,-55.5,100</points>
<connection>
<GID>478</GID>
<name>OUT</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65,91.5,-63.5,91.5</points>
<connection>
<GID>466</GID>
<name>J</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-65,87.5,-63.5,87.5</points>
<connection>
<GID>466</GID>
<name>K</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,87,-48.5,99</points>
<intersection>87 4</intersection>
<intersection>91 2</intersection>
<intersection>99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,99,-40.5,99</points>
<connection>
<GID>479</GID>
<name>OUT</name></connection>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48.5,91,-47.5,91</points>
<connection>
<GID>469</GID>
<name>J</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-48.5,87,-47.5,87</points>
<connection>
<GID>469</GID>
<name>K</name></connection>
<intersection>-48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,87.5,-33,98</points>
<intersection>87.5 4</intersection>
<intersection>91.5 2</intersection>
<intersection>98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,98,-23,98</points>
<connection>
<GID>481</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>-33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,91.5,-31.5,91.5</points>
<connection>
<GID>472</GID>
<name>J</name></connection>
<intersection>-33 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-33,87.5,-31.5,87.5</points>
<connection>
<GID>472</GID>
<name>K</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,87.5,-16,97</points>
<intersection>87.5 4</intersection>
<intersection>91.5 2</intersection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,97,-16,97</points>
<connection>
<GID>482</GID>
<name>OUT</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16,91.5,-14.5,91.5</points>
<connection>
<GID>474</GID>
<name>J</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-16,87.5,-14.5,87.5</points>
<connection>
<GID>474</GID>
<name>K</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,91.5,-79.5,91.5</points>
<connection>
<GID>462</GID>
<name>Q</name></connection>
<connection>
<GID>464</GID>
<name>J</name></connection>
<intersection>-86 3</intersection>
<intersection>-83.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-86,56.5,-86,91.5</points>
<intersection>56.5 10</intersection>
<intersection>72 4</intersection>
<intersection>87.5 9</intersection>
<intersection>91.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-86,72,-4.5,72</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>-86 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-83.5,91.5,-83.5,101</points>
<intersection>91.5 1</intersection>
<intersection>101 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-83.5,101,-72.5,101</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>-83.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-86,87.5,-79.5,87.5</points>
<connection>
<GID>464</GID>
<name>K</name></connection>
<intersection>-86 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-86,56.5,-84,56.5</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>-86 3</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,56.5,-72.5,99</points>
<connection>
<GID>478</GID>
<name>IN_1</name></connection>
<intersection>56.5 8</intersection>
<intersection>73 1</intersection>
<intersection>91.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72.5,73,-4.5,73</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>-72.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-73.5,91.5,-72.5,91.5</points>
<connection>
<GID>464</GID>
<name>Q</name></connection>
<intersection>-72.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-72.5,56.5,-67.5,56.5</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>-72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,75,-4.5,75</points>
<connection>
<GID>475</GID>
<name>IN_3</name></connection>
<intersection>-40.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40.5,56.5,-40.5,101</points>
<connection>
<GID>481</GID>
<name>IN_1</name></connection>
<intersection>56.5 9</intersection>
<intersection>75 1</intersection>
<intersection>91 4</intersection>
<intersection>101 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-41.5,91,-40.5,91</points>
<connection>
<GID>469</GID>
<name>Q</name></connection>
<intersection>-40.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-40.5,101,-1,101</points>
<connection>
<GID>484</GID>
<name>IN_1</name></connection>
<intersection>-40.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-40.5,56.5,-36,56.5</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>-40.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,56.5,-56.5,103</points>
<intersection>56.5 9</intersection>
<intersection>74 4</intersection>
<intersection>91.5 3</intersection>
<intersection>98 2</intersection>
<intersection>103 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-56.5,98,-55.5,98</points>
<connection>
<GID>479</GID>
<name>IN_1</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-57.5,91.5,-56.5,91.5</points>
<connection>
<GID>466</GID>
<name>Q</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-56.5,74,-4.5,74</points>
<connection>
<GID>475</GID>
<name>IN_2</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-56.5,103,-1,103</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-56.5,56.5,-53,56.5</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,56.5,-24.5,99</points>
<intersection>56.5 8</intersection>
<intersection>76 3</intersection>
<intersection>91.5 1</intersection>
<intersection>99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25.5,91.5,-24.5,91.5</points>
<connection>
<GID>472</GID>
<name>Q</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,99,-1,99</points>
<connection>
<GID>484</GID>
<name>IN_2</name></connection>
<intersection>-24.5 0</intersection>
<intersection>-23 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-24.5,76,-4.5,76</points>
<connection>
<GID>475</GID>
<name>IN_4</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-23,96,-23,99</points>
<connection>
<GID>482</GID>
<name>IN_1</name></connection>
<intersection>99 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-24.5,56.5,-20,56.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>-24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,56.5,-6.5,97</points>
<intersection>56.5 5</intersection>
<intersection>77 2</intersection>
<intersection>91.5 1</intersection>
<intersection>97 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,91.5,-6.5,91.5</points>
<connection>
<GID>474</GID>
<name>Q</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,77,-4.5,77</points>
<connection>
<GID>475</GID>
<name>IN_5</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-6.5,97,-1,97</points>
<connection>
<GID>484</GID>
<name>IN_3</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-6.5,56.5,-2,56.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,4.5,424.5,4.5</points>
<intersection>-76.5 3</intersection>
<intersection>424.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-76.5,4.5,-76.5,56.5</points>
<intersection>4.5 1</intersection>
<intersection>42 7</intersection>
<intersection>56.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-78,56.5,-76.5,56.5</points>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection>
<intersection>-76.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>424.5,-1566,424.5,4.5</points>
<intersection>-1566 56</intersection>
<intersection>-1344.5 54</intersection>
<intersection>-1105 53</intersection>
<intersection>-846.5 52</intersection>
<intersection>-680 51</intersection>
<intersection>-498 50</intersection>
<intersection>-349 49</intersection>
<intersection>-222 23</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-76.5,42,16,42</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>-76.5 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>244.5,-222,424.5,-222</points>
<intersection>244.5 29</intersection>
<intersection>424.5 5</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>244.5,-225.5,244.5,-222</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>-222 23</intersection></vsegment>
<hsegment>
<ID>49</ID>
<points>334.5,-349,424.5,-349</points>
<connection>
<GID>2094</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>336,-498,424.5,-498</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>338.5,-680,424.5,-680</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>351,-846.5,424.5,-846.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>342,-1105,424.5,-1105</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>342.5,-1344.5,424.5,-1344.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>360,-1566,424.5,-1566</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>424.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-60,9,421,9</points>
<intersection>-60 3</intersection>
<intersection>421 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-60,9,-60,56.5</points>
<intersection>9 1</intersection>
<intersection>43 7</intersection>
<intersection>56.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-61.5,56.5,-60,56.5</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<intersection>-60 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>421,-1557.5,421,9</points>
<intersection>-1557.5 56</intersection>
<intersection>-1335 54</intersection>
<intersection>-1099 53</intersection>
<intersection>-838 30</intersection>
<intersection>-668 52</intersection>
<intersection>-492.5 51</intersection>
<intersection>-346 50</intersection>
<intersection>-220 19</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-60,43,16,43</points>
<connection>
<GID>493</GID>
<name>IN_1</name></connection>
<intersection>-60 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>258,-220,421,-220</points>
<intersection>258 25</intersection>
<intersection>421 5</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>258,-225.5,258,-220</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>-220 19</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>363,-838,421,-838</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>348,-346,421,-346</points>
<connection>
<GID>2096</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>351.5,-492.5,421,-492.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>348.5,-668,421,-668</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>353,-1099,421,-1099</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment>
<hsegment>
<ID>54</ID>
<points>353.5,-1335,421,-1335</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>372,-1557.5,421,-1557.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>421 5</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,13.5,418.5,13.5</points>
<intersection>-46 3</intersection>
<intersection>418.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-46,13.5,-46,56.5</points>
<intersection>13.5 1</intersection>
<intersection>44 7</intersection>
<intersection>56.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-47,56.5,-46,56.5</points>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection>
<intersection>-46 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>418.5,-1547.5,418.5,13.5</points>
<intersection>-1547.5 52</intersection>
<intersection>-1325.5 50</intersection>
<intersection>-1089.5 49</intersection>
<intersection>-828 48</intersection>
<intersection>-659.5 47</intersection>
<intersection>-484.5 21</intersection>
<intersection>-338.5 46</intersection>
<intersection>-217.5 19</intersection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-46,44,16,44</points>
<connection>
<GID>493</GID>
<name>IN_2</name></connection>
<intersection>-46 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>271,-217.5,418.5,-217.5</points>
<intersection>271 25</intersection>
<intersection>418.5 5</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>352,-484.5,418.5,-484.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>271,-225.5,271,-217.5</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>-217.5 19</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>347.5,-338.5,418.5,-338.5</points>
<connection>
<GID>2098</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>348.5,-659.5,418.5,-659.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>363,-828,418.5,-828</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>353,-1089.5,418.5,-1089.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>353,-1325.5,418.5,-1325.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>373.5,-1547.5,418.5,-1547.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>418.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,18,416.5,18</points>
<intersection>-27.5 3</intersection>
<intersection>416.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,18,-27.5,56.5</points>
<intersection>18 1</intersection>
<intersection>45 7</intersection>
<intersection>56.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-30,56.5,-27.5,56.5</points>
<connection>
<GID>490</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>416.5,-1538,416.5,18</points>
<intersection>-1538 53</intersection>
<intersection>-1317 51</intersection>
<intersection>-1080 50</intersection>
<intersection>-821 49</intersection>
<intersection>-652 48</intersection>
<intersection>-476.5 23</intersection>
<intersection>-330.5 47</intersection>
<intersection>-215 21</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-27.5,45,16,45</points>
<connection>
<GID>493</GID>
<name>IN_3</name></connection>
<intersection>-27.5 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>284,-215,416.5,-215</points>
<intersection>284 27</intersection>
<intersection>416.5 5</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>353,-476.5,416.5,-476.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>284,-225.5,284,-215</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>-215 21</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>348.5,-330.5,416.5,-330.5</points>
<connection>
<GID>2100</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>349.5,-652,416.5,-652</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>364.5,-821,416.5,-821</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>354,-1080,416.5,-1080</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>353.5,-1317,416.5,-1317</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment>
<hsegment>
<ID>53</ID>
<points>374,-1538,416.5,-1538</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>416.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12.5,21,412.5,21</points>
<intersection>-12.5 3</intersection>
<intersection>412.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-12.5,21,-12.5,56.5</points>
<intersection>21 1</intersection>
<intersection>46 7</intersection>
<intersection>56.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-14,56.5,-12.5,56.5</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>412.5,-1529.5,412.5,21</points>
<intersection>-1529.5 49</intersection>
<intersection>-1308.5 47</intersection>
<intersection>-1071.5 46</intersection>
<intersection>-811.5 45</intersection>
<intersection>-643 44</intersection>
<intersection>-466 19</intersection>
<intersection>-324.5 43</intersection>
<intersection>-212 17</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-12.5,46,16,46</points>
<connection>
<GID>493</GID>
<name>IN_4</name></connection>
<intersection>-12.5 3</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>296.5,-212,412.5,-212</points>
<intersection>296.5 23</intersection>
<intersection>412.5 5</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>353.5,-466,412.5,-466</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>296.5,-226,296.5,-212</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>-212 17</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>348.5,-324.5,412.5,-324.5</points>
<connection>
<GID>2102</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>350,-643,412.5,-643</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>365,-811.5,412.5,-811.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>354.5,-1071.5,412.5,-1071.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>353.5,-1308.5,412.5,-1308.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>373.5,-1529.5,412.5,-1529.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>412.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,26,10,56.5</points>
<intersection>26 5</intersection>
<intersection>47 8</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,56.5,10,56.5</points>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>10,26,408,26</points>
<intersection>10 0</intersection>
<intersection>408 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>408,-1521,408,26</points>
<intersection>-1521 50</intersection>
<intersection>-1301 48</intersection>
<intersection>-1063 47</intersection>
<intersection>-804.5 46</intersection>
<intersection>-635 45</intersection>
<intersection>-455 20</intersection>
<intersection>-319 44</intersection>
<intersection>-208 18</intersection>
<intersection>26 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10,47,16,47</points>
<connection>
<GID>493</GID>
<name>IN_5</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>309,-208,408,-208</points>
<intersection>309 24</intersection>
<intersection>408 6</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>353,-455,408,-455</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>309,-226,309,-208</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>-208 18</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>349,-319,408,-319</points>
<connection>
<GID>2104</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>350.5,-635,408,-635</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>365.5,-804.5,408,-804.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>355.5,-1063,408,-1063</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>354,-1301,408,-1301</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>373,-1521,408,-1521</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>408 6</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-96.5,91.5,-96.5,112.5</points>
<intersection>91.5 17</intersection>
<intersection>112.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-235.5,112.5,25,112.5</points>
<intersection>-235.5 11</intersection>
<intersection>-96.5 3</intersection>
<intersection>-93 44</intersection>
<intersection>25 43</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-235.5,164.5,-221.5,164.5</points>
<connection>
<GID>450</GID>
<name>J</name></connection>
<intersection>-235.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-235.5,99,-235.5,164.5</points>
<intersection>99 22</intersection>
<intersection>112 23</intersection>
<intersection>112.5 4</intersection>
<intersection>151 21</intersection>
<intersection>158.5 28</intersection>
<intersection>160.5 14</intersection>
<intersection>164.5 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-235.5,160.5,-221.5,160.5</points>
<connection>
<GID>450</GID>
<name>K</name></connection>
<intersection>-235.5 11</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-96.5,91.5,-93,91.5</points>
<connection>
<GID>462</GID>
<name>J</name></connection>
<intersection>-96.5 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-235.5,151,-234,151</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>-235.5 11</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-238,99,-235.5,99</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<intersection>-235.5 11</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-235.5,112,-227,112</points>
<intersection>-235.5 11</intersection>
<intersection>-227 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-227,107.5,-227,112</points>
<connection>
<GID>452</GID>
<name>IN_1</name></connection>
<intersection>112 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-242,158.5,-235.5,158.5</points>
<connection>
<GID>510</GID>
<name>OUT</name></connection>
<intersection>-235.5 11</intersection></hsegment>
<vsegment>
<ID>43</ID>
<points>25,85.5,25,112.5</points>
<connection>
<GID>431</GID>
<name>J</name></connection>
<intersection>112.5 4</intersection></vsegment>
<vsegment>
<ID>44</ID>
<points>-93,87.5,-93,112.5</points>
<connection>
<GID>462</GID>
<name>K</name></connection>
<intersection>112.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94,53.5,-94,144.5</points>
<intersection>53.5 8</intersection>
<intersection>89.5 1</intersection>
<intersection>144.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94,89.5,-14.5,89.5</points>
<connection>
<GID>462</GID>
<name>clock</name></connection>
<connection>
<GID>464</GID>
<name>clock</name></connection>
<connection>
<GID>466</GID>
<name>clock</name></connection>
<connection>
<GID>472</GID>
<name>clock</name></connection>
<connection>
<GID>474</GID>
<name>clock</name></connection>
<intersection>-94 0</intersection>
<intersection>-47.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-47.5,89,-47.5,89.5</points>
<connection>
<GID>469</GID>
<name>clock</name></connection>
<intersection>89.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-94,53.5,-2,53.5</points>
<connection>
<GID>485</GID>
<name>clock</name></connection>
<connection>
<GID>487</GID>
<name>clock</name></connection>
<connection>
<GID>488</GID>
<name>clock</name></connection>
<connection>
<GID>490</GID>
<name>clock</name></connection>
<connection>
<GID>491</GID>
<name>clock</name></connection>
<connection>
<GID>492</GID>
<name>clock</name></connection>
<intersection>-94 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-94,144.5,-91.5,144.5</points>
<connection>
<GID>494</GID>
<name>OUT_0</name></connection>
<intersection>-94 0</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-1142,291,-1137</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>-1142 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>293,-1148.5,293,-1142</points>
<connection>
<GID>419</GID>
<name>IN_2</name></connection>
<intersection>-1142 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291,-1142,293,-1142</points>
<intersection>291 0</intersection>
<intersection>293 1</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306,-1142.5,306,-1137</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>-1142.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>295,-1148.5,295,-1142.5</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>-1142.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>295,-1142.5,306,-1142.5</points>
<intersection>295 1</intersection>
<intersection>306 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-1143.5,317.5,-1136.5</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-1143.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>297,-1148.5,297,-1143.5</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-1143.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>297,-1143.5,317.5,-1143.5</points>
<intersection>297 1</intersection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,-1142,330.5,-1137</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>-1142 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>329.5,-1147.5,329.5,-1142</points>
<connection>
<GID>525</GID>
<name>IN_1</name></connection>
<intersection>-1142 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>329.5,-1142,330.5,-1142</points>
<intersection>329.5 1</intersection>
<intersection>330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>343.5,-1142,343.5,-1136.5</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<intersection>-1142 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>331.5,-1147.5,331.5,-1142</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>-1142 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>331.5,-1142,343.5,-1142</points>
<intersection>331.5 1</intersection>
<intersection>343.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-1158,294,-1154.5</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>-1158 8</intersection>
<intersection>-1157.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>307,-1170.5,307,-1157.5</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>-1165.5 7</intersection>
<intersection>-1157.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>294,-1157.5,307,-1157.5</points>
<intersection>294 0</intersection>
<intersection>307 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>307,-1165.5,318.5,-1165.5</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>307 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>243.5,-1158,294,-1158</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-405.5,128.5,-291</points>
<connection>
<GID>1820</GID>
<name>OUT</name></connection>
<intersection>-405.5 13</intersection>
<intersection>-345 1</intersection>
<intersection>-336.5 7</intersection>
<intersection>-328 3</intersection>
<intersection>-320 8</intersection>
<intersection>-311.5 5</intersection>
<intersection>-298.5 15</intersection>
<intersection>-293.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-345,151.5,-345</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>128.5,-328,150.5,-328</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>128.5,-311.5,149.5,-311.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>128.5,-336.5,151,-336.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>128.5,-320,150,-320</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>128.5,-293.5,149.5,-293.5</points>
<intersection>128.5 0</intersection>
<intersection>149.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>149.5,-303,149.5,-293.5</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>-293.5 9</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>128.5,-405.5,339,-405.5</points>
<intersection>128.5 0</intersection>
<intersection>339 16</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>128.5,-298.5,329.5,-298.5</points>
<connection>
<GID>2092</GID>
<name>IN_1</name></connection>
<intersection>128.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>339,-405.5,339,-401</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-405.5 13</intersection></vsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,-1157,330.5,-1153.5</points>
<connection>
<GID>525</GID>
<name>OUT</name></connection>
<intersection>-1157 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>309,-1170.5,309,-1157</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-1167.5 6</intersection>
<intersection>-1160 7</intersection>
<intersection>-1157 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>309,-1157,330.5,-1157</points>
<intersection>309 1</intersection>
<intersection>330.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>309,-1167.5,318.5,-1167.5</points>
<connection>
<GID>561</GID>
<name>IN_1</name></connection>
<intersection>309 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>203,-1160,309,-1160</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>309 1</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>182,-1079.5,241,-1079.5</points>
<connection>
<GID>571</GID>
<name>OUT</name></connection>
<connection>
<GID>558</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-1115.5,264,-1079.5</points>
<connection>
<GID>534</GID>
<name>IN_1</name></connection>
<intersection>-1079.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,-1079.5,264,-1079.5</points>
<connection>
<GID>558</GID>
<name>Q</name></connection>
<intersection>264 0</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181.5,-1069.5,228,-1069.5</points>
<connection>
<GID>573</GID>
<name>OUT</name></connection>
<connection>
<GID>559</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-1115.5,277.5,-1069.5</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<intersection>-1069.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234,-1069.5,277.5,-1069.5</points>
<connection>
<GID>559</GID>
<name>Q</name></connection>
<intersection>277.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180,-1058.5,215,-1058.5</points>
<connection>
<GID>574</GID>
<name>OUT</name></connection>
<connection>
<GID>560</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-1115.5,290.5,-1058.5</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>-1058.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221,-1058.5,290.5,-1058.5</points>
<connection>
<GID>560</GID>
<name>Q</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160.5,-189.5,219.5,-189.5</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<connection>
<GID>543</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-225.5,242.5,-189.5</points>
<connection>
<GID>513</GID>
<name>IN_1</name></connection>
<intersection>-189.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-189.5,242.5,-189.5</points>
<connection>
<GID>543</GID>
<name>Q</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160,-179.5,206.5,-179.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<connection>
<GID>546</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,-225.5,256,-179.5</points>
<connection>
<GID>514</GID>
<name>IN_1</name></connection>
<intersection>-179.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-179.5,256,-179.5</points>
<connection>
<GID>546</GID>
<name>Q</name></connection>
<intersection>256 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158.5,-168.5,193.5,-168.5</points>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<connection>
<GID>547</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-225.5,269,-168.5</points>
<connection>
<GID>516</GID>
<name>IN_1</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-168.5,269,-168.5</points>
<connection>
<GID>547</GID>
<name>Q</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158,-159.5,186,-159.5</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<connection>
<GID>548</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-225.5,282,-159.5</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<intersection>-159.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-159.5,282,-159.5</points>
<connection>
<GID>548</GID>
<name>Q</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-152,177.5,-152</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<connection>
<GID>549</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-226,294.5,-152</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-152,294.5,-152</points>
<connection>
<GID>549</GID>
<name>Q</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-144.5,168.5,-144.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<connection>
<GID>550</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307,-226,307,-144.5</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>-144.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174.5,-144.5,307,-144.5</points>
<connection>
<GID>550</GID>
<name>Q</name></connection>
<intersection>307 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,-346,209.5,-346</points>
<connection>
<GID>528</GID>
<name>OUT</name></connection>
<connection>
<GID>551</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-1049.5,207.5,-1049.5</points>
<connection>
<GID>575</GID>
<name>OUT</name></connection>
<connection>
<GID>563</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>303.5,-1115.5,303.5,-1049.5</points>
<connection>
<GID>539</GID>
<name>IN_1</name></connection>
<intersection>-1049.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-1049.5,303.5,-1049.5</points>
<connection>
<GID>563</GID>
<name>Q</name></connection>
<intersection>303.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>178.5,-1042,199,-1042</points>
<connection>
<GID>576</GID>
<name>OUT</name></connection>
<connection>
<GID>565</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-1116,316,-1042</points>
<connection>
<GID>540</GID>
<name>IN_1</name></connection>
<intersection>-1042 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205,-1042,316,-1042</points>
<connection>
<GID>565</GID>
<name>Q</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177.5,-1034.5,190,-1034.5</points>
<connection>
<GID>577</GID>
<name>OUT</name></connection>
<connection>
<GID>567</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-1116,328.5,-1034.5</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>-1034.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196,-1034.5,328.5,-1034.5</points>
<connection>
<GID>567</GID>
<name>Q</name></connection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-1081.5,185,-1030.5</points>
<connection>
<GID>569</GID>
<name>OUT_0</name></connection>
<intersection>-1081.5 7</intersection>
<intersection>-1071.5 5</intersection>
<intersection>-1060.5 8</intersection>
<intersection>-1051.5 3</intersection>
<intersection>-1044 9</intersection>
<intersection>-1036.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-1036.5,190,-1036.5</points>
<connection>
<GID>567</GID>
<name>clock</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185,-1051.5,207.5,-1051.5</points>
<connection>
<GID>563</GID>
<name>clock</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>185,-1071.5,228,-1071.5</points>
<connection>
<GID>559</GID>
<name>clock</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>185,-1081.5,241,-1081.5</points>
<connection>
<GID>558</GID>
<name>clock</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>185,-1060.5,215,-1060.5</points>
<connection>
<GID>560</GID>
<name>clock</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185,-1044,199,-1044</points>
<connection>
<GID>565</GID>
<name>clock</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-1402.5,147,-1247.5</points>
<connection>
<GID>1841</GID>
<name>OUT</name></connection>
<intersection>-1402.5 13</intersection>
<intersection>-1312.5 1</intersection>
<intersection>-1302.5 3</intersection>
<intersection>-1291.5 5</intersection>
<intersection>-1282.5 7</intersection>
<intersection>-1275 9</intersection>
<intersection>-1251 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-1312.5,178,-1312.5</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>147,-1302.5,177.5,-1302.5</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>147,-1291.5,176,-1291.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>147,-1282.5,175.5,-1282.5</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>147,-1275,174.5,-1275</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>147,-1251,332.5,-1251</points>
<intersection>147 0</intersection>
<intersection>173.5 15</intersection>
<intersection>332.5 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>147,-1402.5,332.5,-1402.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>147 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>332.5,-1251,332.5,-1188.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>-1251 11</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>173.5,-1267.5,173.5,-1251</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>-1251 11</intersection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267,-1359,267,-1355.5</points>
<connection>
<GID>595</GID>
<name>OUT</name></connection>
<intersection>-1359 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267,-1359,268,-1359</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>267 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-1359.5,280.5,-1355.5</points>
<connection>
<GID>596</GID>
<name>OUT</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280.5,-1359.5,284,-1359.5</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,-1359.5,293.5,-1355.5</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293.5,-1359.5,297.5,-1359.5</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-1359.5,309.5,-1355.5</points>
<intersection>-1359.5 1</intersection>
<intersection>-1355.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309.5,-1359.5,312.5,-1359.5</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>306.5,-1355.5,309.5,-1355.5</points>
<connection>
<GID>598</GID>
<name>OUT</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-1358,319,-1356</points>
<connection>
<GID>599</GID>
<name>OUT</name></connection>
<intersection>-1358 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-1358,323,-1358</points>
<intersection>319 0</intersection>
<intersection>323 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>323,-1359.5,323,-1358</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>-1358 1</intersection></vsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,-1358,331.5,-1356</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<intersection>-1358 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331.5,-1358,336,-1358</points>
<intersection>331.5 0</intersection>
<intersection>336 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>336,-1359.5,336,-1358</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>-1358 1</intersection></vsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-1367,278,-1359</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>-1359 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-1359,278,-1359</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-1367,293,-1359.5</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-1359.5,293,-1359.5</points>
<connection>
<GID>579</GID>
<name>OUT_0</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-1367,308,-1359.5</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-1359.5,308,-1359.5</points>
<connection>
<GID>580</GID>
<name>OUT_0</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-1366.5,319.5,-1359.5</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-1359.5,319.5,-1359.5</points>
<connection>
<GID>581</GID>
<name>OUT_0</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-1367,332.5,-1359.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>329,-1359.5,332.5,-1359.5</points>
<connection>
<GID>582</GID>
<name>OUT_0</name></connection>
<intersection>332.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345.5,-1366.5,345.5,-1359.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>-1359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-1359.5,345.5,-1359.5</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>345.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-1376.5,278,-1371</points>
<connection>
<GID>584</GID>
<name>OUT_0</name></connection>
<intersection>-1376.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>293,-1382.5,293,-1376.5</points>
<connection>
<GID>591</GID>
<name>IN_3</name></connection>
<intersection>-1376.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>278,-1376.5,293,-1376.5</points>
<intersection>278 0</intersection>
<intersection>293 1</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-1376,293,-1371</points>
<connection>
<GID>585</GID>
<name>OUT_0</name></connection>
<intersection>-1376 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>295,-1382.5,295,-1376</points>
<connection>
<GID>591</GID>
<name>IN_2</name></connection>
<intersection>-1376 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>293,-1376,295,-1376</points>
<intersection>293 0</intersection>
<intersection>295 1</intersection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-1376.5,308,-1371</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>-1376.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>297,-1382.5,297,-1376.5</points>
<connection>
<GID>591</GID>
<name>IN_1</name></connection>
<intersection>-1376.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>297,-1376.5,308,-1376.5</points>
<intersection>297 1</intersection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-1377.5,319.5,-1370.5</points>
<connection>
<GID>587</GID>
<name>OUT_0</name></connection>
<intersection>-1377.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>299,-1382.5,299,-1377.5</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>-1377.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>299,-1377.5,319.5,-1377.5</points>
<intersection>299 1</intersection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-1376,332.5,-1371</points>
<connection>
<GID>588</GID>
<name>OUT_0</name></connection>
<intersection>-1376 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>331.5,-1381.5,331.5,-1376</points>
<connection>
<GID>593</GID>
<name>IN_1</name></connection>
<intersection>-1376 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>331.5,-1376,332.5,-1376</points>
<intersection>331.5 1</intersection>
<intersection>332.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345.5,-1376,345.5,-1370.5</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<intersection>-1376 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>333.5,-1381.5,333.5,-1376</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<intersection>-1376 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>333.5,-1376,345.5,-1376</points>
<intersection>333.5 1</intersection>
<intersection>345.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296,-1391.5,296,-1388.5</points>
<connection>
<GID>591</GID>
<name>OUT</name></connection>
<intersection>-1391.5 2</intersection>
<intersection>-1391.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>309,-1404.5,309,-1391.5</points>
<connection>
<GID>594</GID>
<name>IN_1</name></connection>
<intersection>-1399.5 7</intersection>
<intersection>-1391.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>245.5,-1391.5,309,-1391.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>296 0</intersection>
<intersection>309 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>309,-1399.5,320.5,-1399.5</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>309 1</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332.5,-1391,332.5,-1387.5</points>
<connection>
<GID>593</GID>
<name>OUT</name></connection>
<intersection>-1391 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>311,-1404.5,311,-1391</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>-1401.5 6</intersection>
<intersection>-1393.5 7</intersection>
<intersection>-1391 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>311,-1391,332.5,-1391</points>
<intersection>311 1</intersection>
<intersection>332.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>311,-1401.5,320.5,-1401.5</points>
<connection>
<GID>608</GID>
<name>IN_1</name></connection>
<intersection>311 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>205,-1393.5,311,-1393.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>311 1</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184,-1313.5,243,-1313.5</points>
<connection>
<GID>614</GID>
<name>OUT</name></connection>
<connection>
<GID>605</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-1349.5,266,-1313.5</points>
<connection>
<GID>595</GID>
<name>IN_1</name></connection>
<intersection>-1313.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249,-1313.5,266,-1313.5</points>
<connection>
<GID>605</GID>
<name>Q</name></connection>
<intersection>266 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>183.5,-1303.5,230,-1303.5</points>
<connection>
<GID>615</GID>
<name>OUT</name></connection>
<connection>
<GID>606</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-1349.5,279.5,-1303.5</points>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<intersection>-1303.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-1303.5,279.5,-1303.5</points>
<connection>
<GID>606</GID>
<name>Q</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>182,-1292.5,217,-1292.5</points>
<connection>
<GID>616</GID>
<name>OUT</name></connection>
<connection>
<GID>607</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-1349.5,292.5,-1292.5</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>-1292.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,-1292.5,292.5,-1292.5</points>
<connection>
<GID>607</GID>
<name>Q</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181.5,-1283.5,209.5,-1283.5</points>
<connection>
<GID>617</GID>
<name>OUT</name></connection>
<connection>
<GID>609</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,-1349.5,305.5,-1283.5</points>
<connection>
<GID>598</GID>
<name>IN_1</name></connection>
<intersection>-1283.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-1283.5,305.5,-1283.5</points>
<connection>
<GID>609</GID>
<name>Q</name></connection>
<intersection>305.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180.5,-1276,201,-1276</points>
<connection>
<GID>618</GID>
<name>OUT</name></connection>
<connection>
<GID>610</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318,-1350,318,-1276</points>
<connection>
<GID>599</GID>
<name>IN_1</name></connection>
<intersection>-1276 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-1276,318,-1276</points>
<connection>
<GID>610</GID>
<name>Q</name></connection>
<intersection>318 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-1268.5,192,-1268.5</points>
<connection>
<GID>619</GID>
<name>OUT</name></connection>
<connection>
<GID>611</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,-1350,330.5,-1268.5</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<intersection>-1268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-1268.5,330.5,-1268.5</points>
<connection>
<GID>611</GID>
<name>Q</name></connection>
<intersection>330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-1315.5,187,-1264.5</points>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection>
<intersection>-1315.5 7</intersection>
<intersection>-1305.5 5</intersection>
<intersection>-1294.5 8</intersection>
<intersection>-1285.5 3</intersection>
<intersection>-1278 9</intersection>
<intersection>-1270.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-1270.5,192,-1270.5</points>
<connection>
<GID>611</GID>
<name>clock</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>187,-1285.5,209.5,-1285.5</points>
<connection>
<GID>609</GID>
<name>clock</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>187,-1305.5,230,-1305.5</points>
<connection>
<GID>606</GID>
<name>clock</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>187,-1315.5,243,-1315.5</points>
<connection>
<GID>605</GID>
<name>clock</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>187,-1294.5,217,-1294.5</points>
<connection>
<GID>607</GID>
<name>clock</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>187,-1278,201,-1278</points>
<connection>
<GID>610</GID>
<name>clock</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-1629.5,156,-1461</points>
<intersection>-1629.5 13</intersection>
<intersection>-1539.5 1</intersection>
<intersection>-1529.5 3</intersection>
<intersection>-1518.5 5</intersection>
<intersection>-1509.5 7</intersection>
<intersection>-1502 9</intersection>
<intersection>-1468.5 11</intersection>
<intersection>-1461 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-1539.5,187,-1539.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>156,-1529.5,186.5,-1529.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>156,-1518.5,185,-1518.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>156,-1509.5,184.5,-1509.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>156,-1502,183.5,-1502</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>156,-1468.5,338.5,-1468.5</points>
<intersection>156 0</intersection>
<intersection>182.5 15</intersection>
<intersection>338.5 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>156,-1629.5,341.5,-1629.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>156 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>338.5,-1468.5,338.5,-1426</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>-1468.5 11</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>182.5,-1494.5,182.5,-1468.5</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>-1468.5 11</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>154,-1461,156,-1461</points>
<connection>
<GID>1845</GID>
<name>OUT</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-1586,276,-1582.5</points>
<connection>
<GID>637</GID>
<name>OUT</name></connection>
<intersection>-1586 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-1586,277,-1586</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289.5,-1586.5,289.5,-1582.5</points>
<connection>
<GID>638</GID>
<name>OUT</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289.5,-1586.5,293,-1586.5</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>289.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-1586.5,302.5,-1582.5</points>
<connection>
<GID>639</GID>
<name>OUT</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-1586.5,306.5,-1586.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-1586.5,318.5,-1582.5</points>
<intersection>-1586.5 1</intersection>
<intersection>-1582.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-1586.5,321.5,-1586.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>318.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>315.5,-1582.5,318.5,-1582.5</points>
<connection>
<GID>640</GID>
<name>OUT</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328,-1585,328,-1583</points>
<connection>
<GID>641</GID>
<name>OUT</name></connection>
<intersection>-1585 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>328,-1585,332,-1585</points>
<intersection>328 0</intersection>
<intersection>332 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>332,-1586.5,332,-1585</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>-1585 1</intersection></vsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>340.5,-1585,340.5,-1583</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<intersection>-1585 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>340.5,-1585,345,-1585</points>
<intersection>340.5 0</intersection>
<intersection>345 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>345,-1586.5,345,-1585</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>-1585 1</intersection></vsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-1594,287,-1586</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-1586 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283,-1586,287,-1586</points>
<connection>
<GID>662</GID>
<name>OUT_0</name></connection>
<intersection>287 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-1594,302,-1586.5</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>299,-1586.5,302,-1586.5</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<intersection>302 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-1594,317,-1586.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-1586.5,317,-1586.5</points>
<connection>
<GID>622</GID>
<name>OUT_0</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-1593.5,328.5,-1586.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,-1586.5,328.5,-1586.5</points>
<connection>
<GID>623</GID>
<name>OUT_0</name></connection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-1594,341.5,-1586.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>338,-1586.5,341.5,-1586.5</points>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<intersection>341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-1593.5,354.5,-1586.5</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>-1586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,-1586.5,354.5,-1586.5</points>
<connection>
<GID>625</GID>
<name>OUT_0</name></connection>
<intersection>354.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-1603.5,287,-1598</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<intersection>-1603.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>302,-1609.5,302,-1603.5</points>
<connection>
<GID>633</GID>
<name>IN_3</name></connection>
<intersection>-1603.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>287,-1603.5,302,-1603.5</points>
<intersection>287 0</intersection>
<intersection>302 1</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-1603,302,-1598</points>
<connection>
<GID>627</GID>
<name>OUT_0</name></connection>
<intersection>-1603 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>304,-1609.5,304,-1603</points>
<connection>
<GID>633</GID>
<name>IN_2</name></connection>
<intersection>-1603 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>302,-1603,304,-1603</points>
<intersection>302 0</intersection>
<intersection>304 1</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-1603.5,317,-1598</points>
<connection>
<GID>628</GID>
<name>OUT_0</name></connection>
<intersection>-1603.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>306,-1609.5,306,-1603.5</points>
<connection>
<GID>633</GID>
<name>IN_1</name></connection>
<intersection>-1603.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>306,-1603.5,317,-1603.5</points>
<intersection>306 1</intersection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,-1604.5,328.5,-1597.5</points>
<connection>
<GID>629</GID>
<name>OUT_0</name></connection>
<intersection>-1604.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>308,-1609.5,308,-1604.5</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-1604.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>308,-1604.5,328.5,-1604.5</points>
<intersection>308 1</intersection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-1603,341.5,-1598</points>
<connection>
<GID>630</GID>
<name>OUT_0</name></connection>
<intersection>-1603 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>340.5,-1608.5,340.5,-1603</points>
<connection>
<GID>635</GID>
<name>IN_1</name></connection>
<intersection>-1603 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>340.5,-1603,341.5,-1603</points>
<intersection>340.5 1</intersection>
<intersection>341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>354.5,-1603,354.5,-1597.5</points>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection>
<intersection>-1603 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>342.5,-1608.5,342.5,-1603</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>-1603 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>342.5,-1603,354.5,-1603</points>
<intersection>342.5 1</intersection>
<intersection>354.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305,-1620,305,-1615.5</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<intersection>-1620 8</intersection>
<intersection>-1618.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>318,-1631.5,318,-1618.5</points>
<connection>
<GID>636</GID>
<name>IN_1</name></connection>
<intersection>-1626.5 7</intersection>
<intersection>-1618.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>305,-1618.5,318,-1618.5</points>
<intersection>305 0</intersection>
<intersection>318 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>318,-1626.5,329.5,-1626.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>318 1</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>268,-1620,305,-1620</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>305 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341.5,-1618,341.5,-1614.5</points>
<connection>
<GID>635</GID>
<name>OUT</name></connection>
<intersection>-1618 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>320,-1631.5,320,-1618</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>-1628.5 6</intersection>
<intersection>-1622 7</intersection>
<intersection>-1618 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>320,-1618,341.5,-1618</points>
<intersection>320 1</intersection>
<intersection>341.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>320,-1628.5,329.5,-1628.5</points>
<connection>
<GID>650</GID>
<name>IN_1</name></connection>
<intersection>320 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>227.5,-1622,320,-1622</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>320 1</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>193,-1540.5,252,-1540.5</points>
<connection>
<GID>656</GID>
<name>OUT</name></connection>
<connection>
<GID>647</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-1576.5,275,-1540.5</points>
<connection>
<GID>637</GID>
<name>IN_1</name></connection>
<intersection>-1540.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,-1540.5,275,-1540.5</points>
<connection>
<GID>647</GID>
<name>Q</name></connection>
<intersection>275 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192.5,-1530.5,239,-1530.5</points>
<connection>
<GID>657</GID>
<name>OUT</name></connection>
<connection>
<GID>648</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-1576.5,288.5,-1530.5</points>
<connection>
<GID>638</GID>
<name>IN_1</name></connection>
<intersection>-1530.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-1530.5,288.5,-1530.5</points>
<connection>
<GID>648</GID>
<name>Q</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191,-1519.5,226,-1519.5</points>
<connection>
<GID>658</GID>
<name>OUT</name></connection>
<connection>
<GID>649</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-1576.5,301.5,-1519.5</points>
<connection>
<GID>639</GID>
<name>IN_1</name></connection>
<intersection>-1519.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232,-1519.5,301.5,-1519.5</points>
<connection>
<GID>649</GID>
<name>Q</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190.5,-1510.5,218.5,-1510.5</points>
<connection>
<GID>659</GID>
<name>OUT</name></connection>
<connection>
<GID>651</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314.5,-1576.5,314.5,-1510.5</points>
<connection>
<GID>640</GID>
<name>IN_1</name></connection>
<intersection>-1510.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224.5,-1510.5,314.5,-1510.5</points>
<connection>
<GID>651</GID>
<name>Q</name></connection>
<intersection>314.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,-1503,210,-1503</points>
<connection>
<GID>660</GID>
<name>OUT</name></connection>
<connection>
<GID>652</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327,-1577,327,-1503</points>
<connection>
<GID>641</GID>
<name>IN_1</name></connection>
<intersection>-1503 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,-1503,327,-1503</points>
<connection>
<GID>652</GID>
<name>Q</name></connection>
<intersection>327 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,-1495.5,201,-1495.5</points>
<connection>
<GID>661</GID>
<name>OUT</name></connection>
<connection>
<GID>653</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,-1577,339.5,-1495.5</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>-1495.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-1495.5,339.5,-1495.5</points>
<connection>
<GID>653</GID>
<name>Q</name></connection>
<intersection>339.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-1542.5,196,-1491.5</points>
<connection>
<GID>654</GID>
<name>OUT_0</name></connection>
<intersection>-1542.5 7</intersection>
<intersection>-1532.5 5</intersection>
<intersection>-1521.5 8</intersection>
<intersection>-1512.5 3</intersection>
<intersection>-1505 9</intersection>
<intersection>-1497.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196,-1497.5,201,-1497.5</points>
<connection>
<GID>653</GID>
<name>clock</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>196,-1512.5,218.5,-1512.5</points>
<connection>
<GID>651</GID>
<name>clock</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>196,-1532.5,239,-1532.5</points>
<connection>
<GID>648</GID>
<name>clock</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>196,-1542.5,252,-1542.5</points>
<connection>
<GID>647</GID>
<name>clock</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>196,-1521.5,226,-1521.5</points>
<connection>
<GID>649</GID>
<name>clock</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>196,-1505,210,-1505</points>
<connection>
<GID>652</GID>
<name>clock</name></connection>
<intersection>196 0</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-350.5,242,-346</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>-346 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-346,242,-346</points>
<connection>
<GID>551</GID>
<name>Q</name></connection>
<intersection>242 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-337.5,201.5,-337.5</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<connection>
<GID>552</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-350.5,255.5,-337.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>-337.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-337.5,255.5,-337.5</points>
<connection>
<GID>552</GID>
<name>Q</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-329,194.5,-329</points>
<connection>
<GID>530</GID>
<name>OUT</name></connection>
<connection>
<GID>553</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-350.5,268.5,-329</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<intersection>-329 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,-329,268.5,-329</points>
<connection>
<GID>553</GID>
<name>Q</name></connection>
<intersection>268.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,-321,185.5,-321</points>
<connection>
<GID>531</GID>
<name>OUT</name></connection>
<connection>
<GID>554</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-350.5,281.5,-321</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>-321 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-321,281.5,-321</points>
<connection>
<GID>554</GID>
<name>Q</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-133,122.5,-132.5</points>
<connection>
<GID>1818</GID>
<name>IN_1</name></connection>
<intersection>-132.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>119,-132.5,119,-128.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>119,-132.5,122.5,-132.5</points>
<intersection>119 1</intersection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155.5,-312.5,178.5,-312.5</points>
<connection>
<GID>532</GID>
<name>OUT</name></connection>
<connection>
<GID>555</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-133,124.5,-132.5</points>
<connection>
<GID>1818</GID>
<name>IN_0</name></connection>
<intersection>-132.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>131,-132.5,131,-128</points>
<connection>
<GID>1814</GID>
<name>OUT_0</name></connection>
<intersection>-132.5 2</intersection>
<intersection>-128 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-132.5,131,-132.5</points>
<intersection>124.5 0</intersection>
<intersection>131 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>131,-128,153,-128</points>
<intersection>131 1</intersection>
<intersection>153 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>153,-128,153,-126</points>
<connection>
<GID>1850</GID>
<name>N_in0</name></connection>
<intersection>-128 4</intersection></vsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-351,294,-312.5</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>-312.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-312.5,294,-312.5</points>
<connection>
<GID>555</GID>
<name>Q</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>2141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-285,123.5,-281.5</points>
<connection>
<GID>526</GID>
<name>OUT_0</name></connection>
<intersection>-285 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>123.5,-285,127.5,-285</points>
<connection>
<GID>1820</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155.5,-304,170.5,-304</points>
<connection>
<GID>533</GID>
<name>OUT</name></connection>
<connection>
<GID>556</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>2142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-285,129.5,-283</points>
<connection>
<GID>1820</GID>
<name>IN_0</name></connection>
<intersection>-283 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>130,-283,130,-281.5</points>
<connection>
<GID>1822</GID>
<name>OUT_0</name></connection>
<intersection>-283 2</intersection>
<intersection>-282.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-283,130,-283</points>
<intersection>129.5 0</intersection>
<intersection>130 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130,-282.5,141,-282.5</points>
<intersection>130 1</intersection>
<intersection>141 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>141,-282.5,141,-280.5</points>
<connection>
<GID>1853</GID>
<name>N_in0</name></connection>
<intersection>-282.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306.5,-351,306.5,-304</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>-304 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176.5,-304,306.5,-304</points>
<connection>
<GID>556</GID>
<name>Q</name></connection>
<intersection>306.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-408.5,114.5,-405</points>
<connection>
<GID>1828</GID>
<name>OUT_0</name></connection>
<intersection>-408.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>114.5,-408.5,118.5,-408.5</points>
<connection>
<GID>1825</GID>
<name>IN_1</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-408.5,120.5,-406.5</points>
<connection>
<GID>1825</GID>
<name>IN_0</name></connection>
<intersection>-406.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>121,-406.5,121,-405</points>
<connection>
<GID>1826</GID>
<name>OUT_0</name></connection>
<intersection>-406.5 2</intersection>
<intersection>-405.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120.5,-406.5,121,-406.5</points>
<intersection>120.5 0</intersection>
<intersection>121 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>121,-405.5,131.5,-405.5</points>
<intersection>121 1</intersection>
<intersection>131.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>131.5,-405.5,131.5,-403.5</points>
<connection>
<GID>1854</GID>
<name>N_in0</name></connection>
<intersection>-405.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>2145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-584.5,129,-581</points>
<connection>
<GID>1832</GID>
<name>OUT_0</name></connection>
<intersection>-584.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>129,-584.5,132,-584.5</points>
<intersection>129 0</intersection>
<intersection>132 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>132,-585,132,-584.5</points>
<connection>
<GID>1829</GID>
<name>IN_1</name></connection>
<intersection>-584.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>2146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-585,134,-582.5</points>
<connection>
<GID>1829</GID>
<name>IN_0</name></connection>
<intersection>-582.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>136,-582.5,136,-581</points>
<connection>
<GID>1830</GID>
<name>OUT_0</name></connection>
<intersection>-582.5 2</intersection>
<intersection>-581 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134,-582.5,136,-582.5</points>
<intersection>134 0</intersection>
<intersection>136 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136,-581,147.5,-581</points>
<connection>
<GID>1855</GID>
<name>N_in0</name></connection>
<intersection>136 1</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-348,165.5,-296</points>
<connection>
<GID>566</GID>
<name>OUT_0</name></connection>
<intersection>-348 7</intersection>
<intersection>-339.5 5</intersection>
<intersection>-331 8</intersection>
<intersection>-323 3</intersection>
<intersection>-314.5 9</intersection>
<intersection>-306 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165.5,-306,170.5,-306</points>
<connection>
<GID>556</GID>
<name>clock</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>165.5,-323,185.5,-323</points>
<connection>
<GID>554</GID>
<name>clock</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-339.5,201.5,-339.5</points>
<connection>
<GID>552</GID>
<name>clock</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>165.5,-348,209.5,-348</points>
<connection>
<GID>551</GID>
<name>clock</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>165.5,-331,194.5,-331</points>
<connection>
<GID>553</GID>
<name>clock</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>165.5,-314.5,178.5,-314.5</points>
<connection>
<GID>555</GID>
<name>clock</name></connection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-782,147.5,-778.5</points>
<connection>
<GID>1836</GID>
<name>OUT_0</name></connection>
<intersection>-782 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>147.5,-782,151.5,-782</points>
<connection>
<GID>1833</GID>
<name>IN_1</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-191.5,163,-140.5</points>
<connection>
<GID>568</GID>
<name>OUT_0</name></connection>
<intersection>-191.5 7</intersection>
<intersection>-181.5 5</intersection>
<intersection>-170.5 8</intersection>
<intersection>-161.5 3</intersection>
<intersection>-154 9</intersection>
<intersection>-146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-146.5,168.5,-146.5</points>
<connection>
<GID>550</GID>
<name>clock</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>163,-161.5,186,-161.5</points>
<connection>
<GID>548</GID>
<name>clock</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>163,-181.5,206.5,-181.5</points>
<connection>
<GID>546</GID>
<name>clock</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>163,-191.5,219.5,-191.5</points>
<connection>
<GID>543</GID>
<name>clock</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>163,-170.5,193.5,-170.5</points>
<connection>
<GID>547</GID>
<name>clock</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>163,-154,177.5,-154</points>
<connection>
<GID>549</GID>
<name>clock</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>2148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-782,153.5,-780</points>
<connection>
<GID>1833</GID>
<name>IN_0</name></connection>
<intersection>-780 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>154,-780,154,-778.5</points>
<connection>
<GID>1834</GID>
<name>OUT_0</name></connection>
<intersection>-780 2</intersection>
<intersection>-779 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>153.5,-780,154,-780</points>
<intersection>153.5 0</intersection>
<intersection>154 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>154,-779,164.5,-779</points>
<connection>
<GID>1856</GID>
<name>N_in0</name></connection>
<intersection>154 1</intersection></hsegment></shape></wire>
<wire>
<ID>2149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-999.5,141,-996</points>
<connection>
<GID>1840</GID>
<name>OUT_0</name></connection>
<intersection>-999.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>141,-999.5,145,-999.5</points>
<connection>
<GID>1837</GID>
<name>IN_1</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388.5,-357.5,388.5,-123</points>
<intersection>-357.5 17</intersection>
<intersection>-195.5 3</intersection>
<intersection>-123 26</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>171.5,-195.5,388.5,-195.5</points>
<connection>
<GID>543</GID>
<name>clear</name></connection>
<intersection>171.5 27</intersection>
<intersection>180.5 28</intersection>
<intersection>189 29</intersection>
<intersection>196.5 30</intersection>
<intersection>209.5 31</intersection>
<intersection>388.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>173.5,-357.5,388.5,-357.5</points>
<intersection>173.5 33</intersection>
<intersection>181.5 34</intersection>
<intersection>188.5 35</intersection>
<intersection>197.5 36</intersection>
<intersection>204.5 37</intersection>
<intersection>212.5 38</intersection>
<intersection>388 39</intersection>
<intersection>388.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>326,-123,388.5,-123</points>
<intersection>326 32</intersection>
<intersection>388.5 0</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>171.5,-195.5,171.5,-150.5</points>
<connection>
<GID>550</GID>
<name>clear</name></connection>
<intersection>-195.5 3</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>180.5,-195.5,180.5,-158</points>
<connection>
<GID>549</GID>
<name>clear</name></connection>
<intersection>-195.5 3</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>189,-195.5,189,-165.5</points>
<connection>
<GID>548</GID>
<name>clear</name></connection>
<intersection>-195.5 3</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>196.5,-195.5,196.5,-174.5</points>
<connection>
<GID>547</GID>
<name>clear</name></connection>
<intersection>-195.5 3</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>209.5,-195.5,209.5,-185.5</points>
<connection>
<GID>546</GID>
<name>clear</name></connection>
<intersection>-195.5 3</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>326,-123,326,-116.5</points>
<connection>
<GID>572</GID>
<name>OUT_0</name></connection>
<intersection>-123 26</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>173.5,-357.5,173.5,-310</points>
<connection>
<GID>556</GID>
<name>clear</name></connection>
<intersection>-357.5 17</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>181.5,-357.5,181.5,-318.5</points>
<connection>
<GID>555</GID>
<name>clear</name></connection>
<intersection>-357.5 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>188.5,-357.5,188.5,-327</points>
<connection>
<GID>554</GID>
<name>clear</name></connection>
<intersection>-357.5 17</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>197.5,-357.5,197.5,-335</points>
<connection>
<GID>553</GID>
<name>clear</name></connection>
<intersection>-357.5 17</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>204.5,-357.5,204.5,-343.5</points>
<connection>
<GID>552</GID>
<name>clear</name></connection>
<intersection>-357.5 17</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>212.5,-357.5,212.5,-352</points>
<connection>
<GID>551</GID>
<name>clear</name></connection>
<intersection>-357.5 17</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>388,-1085.5,388,-357.5</points>
<intersection>-1085.5 105</intersection>
<intersection>-863.5 84</intersection>
<intersection>-672 64</intersection>
<intersection>-488.5 43</intersection>
<intersection>-357.5 17</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>180.5,-488.5,388,-488.5</points>
<intersection>180.5 53</intersection>
<intersection>190 54</intersection>
<intersection>198.5 55</intersection>
<intersection>206 56</intersection>
<intersection>219 57</intersection>
<intersection>232 59</intersection>
<intersection>388 39</intersection></hsegment>
<vsegment>
<ID>53</ID>
<points>180.5,-488.5,180.5,-437.5</points>
<intersection>-488.5 43</intersection>
<intersection>-437.5 58</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>190,-488.5,190,-445</points>
<connection>
<GID>130</GID>
<name>clear</name></connection>
<intersection>-488.5 43</intersection></vsegment>
<vsegment>
<ID>55</ID>
<points>198.5,-488.5,198.5,-452.5</points>
<connection>
<GID>129</GID>
<name>clear</name></connection>
<intersection>-488.5 43</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>206,-488.5,206,-461.5</points>
<connection>
<GID>126</GID>
<name>clear</name></connection>
<intersection>-488.5 43</intersection></vsegment>
<vsegment>
<ID>57</ID>
<points>219,-488.5,219,-472.5</points>
<connection>
<GID>125</GID>
<name>clear</name></connection>
<intersection>-488.5 43</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>180.5,-437.5,181,-437.5</points>
<connection>
<GID>134</GID>
<name>clear</name></connection>
<intersection>180.5 53</intersection></hsegment>
<vsegment>
<ID>59</ID>
<points>232,-488.5,232,-482.5</points>
<connection>
<GID>123</GID>
<name>clear</name></connection>
<intersection>-488.5 43</intersection></vsegment>
<hsegment>
<ID>64</ID>
<points>189,-672,388,-672</points>
<intersection>189 74</intersection>
<intersection>198 75</intersection>
<intersection>206.5 76</intersection>
<intersection>214 77</intersection>
<intersection>227 78</intersection>
<intersection>240 79</intersection>
<intersection>388 39</intersection></hsegment>
<vsegment>
<ID>74</ID>
<points>189,-672,189,-619.5</points>
<connection>
<GID>228</GID>
<name>clear</name></connection>
<intersection>-672 64</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>198,-672,198,-627</points>
<connection>
<GID>227</GID>
<name>clear</name></connection>
<intersection>-672 64</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>206.5,-672,206.5,-634.5</points>
<connection>
<GID>226</GID>
<name>clear</name></connection>
<intersection>-672 64</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>214,-672,214,-643.5</points>
<connection>
<GID>224</GID>
<name>clear</name></connection>
<intersection>-672 64</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>227,-672,227,-654.5</points>
<connection>
<GID>223</GID>
<name>clear</name></connection>
<intersection>-672 64</intersection></vsegment>
<vsegment>
<ID>79</ID>
<points>240,-672,240,-664.5</points>
<connection>
<GID>222</GID>
<name>clear</name></connection>
<intersection>-672 64</intersection></vsegment>
<hsegment>
<ID>84</ID>
<points>199.5,-863.5,388,-863.5</points>
<connection>
<GID>305</GID>
<name>clear</name></connection>
<intersection>199.5 94</intersection>
<intersection>208.5 95</intersection>
<intersection>217 100</intersection>
<intersection>224.5 97</intersection>
<intersection>237.5 98</intersection>
<intersection>388 39</intersection></hsegment>
<vsegment>
<ID>94</ID>
<points>199.5,-863.5,199.5,-818.5</points>
<connection>
<GID>311</GID>
<name>clear</name></connection>
<intersection>-863.5 84</intersection></vsegment>
<vsegment>
<ID>95</ID>
<points>208.5,-863.5,208.5,-826</points>
<connection>
<GID>310</GID>
<name>clear</name></connection>
<intersection>-863.5 84</intersection></vsegment>
<vsegment>
<ID>97</ID>
<points>224.5,-863.5,224.5,-842.5</points>
<connection>
<GID>307</GID>
<name>clear</name></connection>
<intersection>-863.5 84</intersection></vsegment>
<vsegment>
<ID>98</ID>
<points>237.5,-863.5,237.5,-853.5</points>
<connection>
<GID>306</GID>
<name>clear</name></connection>
<intersection>-863.5 84</intersection></vsegment>
<vsegment>
<ID>100</ID>
<points>217,-863.5,217,-833.5</points>
<connection>
<GID>309</GID>
<name>clear</name></connection>
<intersection>-863.5 84</intersection></vsegment>
<hsegment>
<ID>105</ID>
<points>193,-1085.5,388,-1085.5</points>
<connection>
<GID>558</GID>
<name>clear</name></connection>
<intersection>193 115</intersection>
<intersection>202 116</intersection>
<intersection>210.5 117</intersection>
<intersection>218 118</intersection>
<intersection>231 119</intersection>
<intersection>387.5 120</intersection>
<intersection>388 39</intersection></hsegment>
<vsegment>
<ID>115</ID>
<points>193,-1085.5,193,-1040.5</points>
<connection>
<GID>567</GID>
<name>clear</name></connection>
<intersection>-1085.5 105</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>202,-1085.5,202,-1048</points>
<connection>
<GID>565</GID>
<name>clear</name></connection>
<intersection>-1085.5 105</intersection></vsegment>
<vsegment>
<ID>117</ID>
<points>210.5,-1085.5,210.5,-1055.5</points>
<connection>
<GID>563</GID>
<name>clear</name></connection>
<intersection>-1085.5 105</intersection></vsegment>
<vsegment>
<ID>118</ID>
<points>218,-1085.5,218,-1064.5</points>
<connection>
<GID>560</GID>
<name>clear</name></connection>
<intersection>-1085.5 105</intersection></vsegment>
<vsegment>
<ID>119</ID>
<points>231,-1085.5,231,-1075.5</points>
<connection>
<GID>559</GID>
<name>clear</name></connection>
<intersection>-1085.5 105</intersection></vsegment>
<vsegment>
<ID>120</ID>
<points>387.5,-1319.5,387.5,-1085.5</points>
<intersection>-1319.5 124</intersection>
<intersection>-1085.5 105</intersection></vsegment>
<hsegment>
<ID>124</ID>
<points>195,-1319.5,387.5,-1319.5</points>
<connection>
<GID>605</GID>
<name>clear</name></connection>
<intersection>195 134</intersection>
<intersection>204 135</intersection>
<intersection>212.5 136</intersection>
<intersection>220 137</intersection>
<intersection>233 138</intersection>
<intersection>387 139</intersection>
<intersection>387.5 120</intersection></hsegment>
<vsegment>
<ID>134</ID>
<points>195,-1319.5,195,-1274.5</points>
<connection>
<GID>611</GID>
<name>clear</name></connection>
<intersection>-1319.5 124</intersection></vsegment>
<vsegment>
<ID>135</ID>
<points>204,-1319.5,204,-1282</points>
<connection>
<GID>610</GID>
<name>clear</name></connection>
<intersection>-1319.5 124</intersection></vsegment>
<vsegment>
<ID>136</ID>
<points>212.5,-1319.5,212.5,-1289.5</points>
<connection>
<GID>609</GID>
<name>clear</name></connection>
<intersection>-1319.5 124</intersection></vsegment>
<vsegment>
<ID>137</ID>
<points>220,-1319.5,220,-1298.5</points>
<connection>
<GID>607</GID>
<name>clear</name></connection>
<intersection>-1319.5 124</intersection></vsegment>
<vsegment>
<ID>138</ID>
<points>233,-1319.5,233,-1309.5</points>
<connection>
<GID>606</GID>
<name>clear</name></connection>
<intersection>-1319.5 124</intersection></vsegment>
<vsegment>
<ID>139</ID>
<points>387,-1546.5,387,-1319.5</points>
<intersection>-1546.5 143</intersection>
<intersection>-1319.5 124</intersection></vsegment>
<hsegment>
<ID>143</ID>
<points>204,-1546.5,387,-1546.5</points>
<connection>
<GID>647</GID>
<name>clear</name></connection>
<intersection>204 154</intersection>
<intersection>213 155</intersection>
<intersection>221.5 156</intersection>
<intersection>229 157</intersection>
<intersection>242 158</intersection>
<intersection>387 139</intersection></hsegment>
<vsegment>
<ID>154</ID>
<points>204,-1546.5,204,-1501.5</points>
<connection>
<GID>653</GID>
<name>clear</name></connection>
<intersection>-1546.5 143</intersection></vsegment>
<vsegment>
<ID>155</ID>
<points>213,-1546.5,213,-1509</points>
<connection>
<GID>652</GID>
<name>clear</name></connection>
<intersection>-1546.5 143</intersection></vsegment>
<vsegment>
<ID>156</ID>
<points>221.5,-1546.5,221.5,-1516.5</points>
<connection>
<GID>651</GID>
<name>clear</name></connection>
<intersection>-1546.5 143</intersection></vsegment>
<vsegment>
<ID>157</ID>
<points>229,-1546.5,229,-1525.5</points>
<connection>
<GID>649</GID>
<name>clear</name></connection>
<intersection>-1546.5 143</intersection></vsegment>
<vsegment>
<ID>158</ID>
<points>242,-1546.5,242,-1536.5</points>
<connection>
<GID>648</GID>
<name>clear</name></connection>
<intersection>-1546.5 143</intersection></vsegment></shape></wire>
<wire>
<ID>2150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-999.5,147,-997.5</points>
<connection>
<GID>1837</GID>
<name>IN_0</name></connection>
<intersection>-997.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>147.5,-997.5,147.5,-996</points>
<connection>
<GID>1838</GID>
<name>OUT_0</name></connection>
<intersection>-997.5 2</intersection>
<intersection>-997.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>147,-997.5,157,-997.5</points>
<connection>
<GID>1857</GID>
<name>N_in0</name></connection>
<intersection>147 0</intersection>
<intersection>147.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-1241.5,142,-1238</points>
<connection>
<GID>1844</GID>
<name>OUT_0</name></connection>
<intersection>-1241.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>142,-1241.5,146,-1241.5</points>
<connection>
<GID>1841</GID>
<name>IN_1</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>2152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-1241.5,148,-1239.5</points>
<connection>
<GID>1841</GID>
<name>IN_0</name></connection>
<intersection>-1239.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>148.5,-1239.5,148.5,-1238</points>
<connection>
<GID>1842</GID>
<name>OUT_0</name></connection>
<intersection>-1239.5 2</intersection>
<intersection>-1238.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148,-1239.5,148.5,-1239.5</points>
<intersection>148 0</intersection>
<intersection>148.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148.5,-1238.5,158.5,-1238.5</points>
<connection>
<GID>1858</GID>
<name>N_in0</name></connection>
<intersection>148.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-1455,149,-1451.5</points>
<connection>
<GID>1848</GID>
<name>OUT_0</name></connection>
<intersection>-1455 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>149,-1455,153,-1455</points>
<connection>
<GID>1845</GID>
<name>IN_1</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>2154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-1455,155,-1453</points>
<connection>
<GID>1845</GID>
<name>IN_0</name></connection>
<intersection>-1453 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>155.5,-1453,155.5,-1451.5</points>
<connection>
<GID>1846</GID>
<name>OUT_0</name></connection>
<intersection>-1453 2</intersection>
<intersection>-1452.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>155,-1453,155.5,-1453</points>
<intersection>155 0</intersection>
<intersection>155.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>155.5,-1452.5,164.5,-1452.5</points>
<connection>
<GID>1859</GID>
<name>N_in0</name></connection>
<intersection>155.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,-283,330.5,-282.5</points>
<intersection>-283 1</intersection>
<intersection>-282.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326,-283,330.5,-283</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>330.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330.5,-282.5,335,-282.5</points>
<connection>
<GID>1611</GID>
<name>IN_0</name></connection>
<intersection>330.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286.5,-288.5,455,-288.5</points>
<intersection>286.5 12</intersection>
<intersection>311.5 5</intersection>
<intersection>335 2</intersection>
<intersection>455 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>335,-288.5,335,-284.5</points>
<connection>
<GID>1611</GID>
<name>IN_1</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>455,-288.5,455,-271.5</points>
<connection>
<GID>1613</GID>
<name>IN_1</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>311.5,-291,311.5,-288.5</points>
<connection>
<GID>2090</GID>
<name>J</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>286.5,-288.5,286.5,-286.5</points>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453,-280,453,-271.5</points>
<connection>
<GID>1613</GID>
<name>IN_0</name></connection>
<intersection>-280 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>341,-280,453,-280</points>
<intersection>341 7</intersection>
<intersection>350 2</intersection>
<intersection>453 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>350,-283,350,-280</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>-280 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>341,-283.5,341,-280</points>
<connection>
<GID>1611</GID>
<name>OUT</name></connection>
<intersection>-280 1</intersection></vsegment></shape></wire>
<wire>
<ID>1414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,89.5,28,102.5</points>
<intersection>89.5 1</intersection>
<intersection>102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,89.5,28,89.5</points>
<connection>
<GID>431</GID>
<name>K</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,102.5,28,102.5</points>
<connection>
<GID>443</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-6.54961,518.319,380.732,326.893</PageViewport>
<gate>
<ID>1544</ID>
<type>CC_PULSE</type>
<position>366,160</position>
<output>
<ID>OUT_0</ID>1384 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>1545</ID>
<type>AA_TOGGLE</type>
<position>432,160</position>
<output>
<ID>OUT_0</ID>1385 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1546</ID>
<type>AA_AND2</type>
<position>359.5,109</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1267 </input>
<output>
<ID>OUT</ID>1372 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1547</ID>
<type>AA_AND2</type>
<position>359,119</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1285 </input>
<output>
<ID>OUT</ID>1374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1548</ID>
<type>AA_AND2</type>
<position>357.5,130</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1286 </input>
<output>
<ID>OUT</ID>1376 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1549</ID>
<type>AA_AND2</type>
<position>357,139</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1287 </input>
<output>
<ID>OUT</ID>1378 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1550</ID>
<type>AA_AND2</type>
<position>356,146.5</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1288 </input>
<output>
<ID>OUT</ID>1380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1551</ID>
<type>AA_AND2</type>
<position>355,154</position>
<input>
<ID>IN_0</ID>1229 </input>
<input>
<ID>IN_1</ID>1289 </input>
<output>
<ID>OUT</ID>1382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1552</ID>
<type>AA_LABEL</type>
<position>68.5,151</position>
<gparam>LABEL_TEXT Checking condition for 60</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1553</ID>
<type>AA_TOGGLE</type>
<position>-61.5,290</position>
<output>
<ID>OUT_0</ID>1254 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1554</ID>
<type>AA_LABEL</type>
<position>270,232</position>
<gparam>LABEL_TEXT Problematic Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1555</ID>
<type>BA_NAND4</type>
<position>247,287</position>
<input>
<ID>IN_0</ID>1271 </input>
<input>
<ID>IN_1</ID>1275 </input>
<input>
<ID>IN_2</ID>1279 </input>
<input>
<ID>IN_3</ID>1284 </input>
<output>
<ID>OUT</ID>1261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1556</ID>
<type>AE_DFF_LOW</type>
<position>48,217</position>
<input>
<ID>IN_0</ID>1262 </input>
<output>
<ID>OUT_0</ID>1267 </output>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1557</ID>
<type>BE_JKFF_LOW_NT</type>
<position>30,261.5</position>
<input>
<ID>J</ID>1290 </input>
<input>
<ID>K</ID>1292 </input>
<output>
<ID>Q</ID>1262 </output>
<input>
<ID>clear</ID>1261 </input>
<input>
<ID>clock</ID>1283 </input>
<output>
<ID>nQ</ID>1263 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1558</ID>
<type>BE_JKFF_LOW_NT</type>
<position>79.5,261</position>
<input>
<ID>J</ID>1302 </input>
<input>
<ID>K</ID>1303 </input>
<output>
<ID>Q</ID>1266 </output>
<input>
<ID>clear</ID>1261 </input>
<input>
<ID>clock</ID>1283 </input>
<output>
<ID>nQ</ID>1269 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1559</ID>
<type>AE_DFF_LOW</type>
<position>91,217.5</position>
<input>
<ID>IN_0</ID>1266 </input>
<output>
<ID>OUT_0</ID>1285 </output>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1560</ID>
<type>BE_JKFF_LOW_NT</type>
<position>105.5,261.5</position>
<input>
<ID>J</ID>1304 </input>
<input>
<ID>K</ID>1305 </input>
<output>
<ID>Q</ID>1271 </output>
<input>
<ID>clear</ID>1261 </input>
<input>
<ID>clock</ID>1283 </input>
<output>
<ID>nQ</ID>1274 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1561</ID>
<type>BE_JKFF_LOW_NT</type>
<position>135.5,261</position>
<input>
<ID>J</ID>1306 </input>
<input>
<ID>K</ID>1307 </input>
<output>
<ID>Q</ID>1275 </output>
<input>
<ID>clear</ID>1261 </input>
<input>
<ID>clock</ID>1283 </input>
<output>
<ID>nQ</ID>1276 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1562</ID>
<type>BE_JKFF_LOW_NT</type>
<position>174,259</position>
<input>
<ID>J</ID>1308 </input>
<input>
<ID>K</ID>1309 </input>
<output>
<ID>Q</ID>1279 </output>
<input>
<ID>clear</ID>1261 </input>
<input>
<ID>clock</ID>1283 </input>
<output>
<ID>nQ</ID>1280 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1563</ID>
<type>BE_JKFF_LOW_NT</type>
<position>222.5,258.5</position>
<input>
<ID>J</ID>1310 </input>
<input>
<ID>K</ID>1311 </input>
<output>
<ID>Q</ID>1284 </output>
<input>
<ID>clear</ID>1261 </input>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1564</ID>
<type>AE_DFF_LOW</type>
<position>120.5,217.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<output>
<ID>OUT_0</ID>1286 </output>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1565</ID>
<type>AA_AND2</type>
<position>46.5,270.5</position>
<input>
<ID>IN_0</ID>1318 </input>
<input>
<ID>IN_1</ID>1262 </input>
<output>
<ID>OUT</ID>1264 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1566</ID>
<type>AE_DFF_LOW</type>
<position>449.5,61.5</position>
<input>
<ID>IN_0</ID>1230 </input>
<output>
<ID>OUT_0</ID>1236 </output>
<input>
<ID>clock</ID>1320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1567</ID>
<type>AA_AND2</type>
<position>45.5,253</position>
<input>
<ID>IN_0</ID>1263 </input>
<input>
<ID>IN_1</ID>1319 </input>
<output>
<ID>OUT</ID>1265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1568</ID>
<type>AA_AND2</type>
<position>87.5,270.5</position>
<input>
<ID>IN_0</ID>1264 </input>
<input>
<ID>IN_1</ID>1266 </input>
<output>
<ID>OUT</ID>1268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1569</ID>
<type>AA_AND2</type>
<position>90,252</position>
<input>
<ID>IN_0</ID>1269 </input>
<input>
<ID>IN_1</ID>1265 </input>
<output>
<ID>OUT</ID>1270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1570</ID>
<type>AA_AND2</type>
<position>117,269</position>
<input>
<ID>IN_0</ID>1268 </input>
<input>
<ID>IN_1</ID>1271 </input>
<output>
<ID>OUT</ID>1272 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1571</ID>
<type>AA_AND2</type>
<position>119.5,250.5</position>
<input>
<ID>IN_0</ID>1274 </input>
<input>
<ID>IN_1</ID>1270 </input>
<output>
<ID>OUT</ID>1273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1572</ID>
<type>AA_AND2</type>
<position>143.5,268</position>
<input>
<ID>IN_0</ID>1272 </input>
<input>
<ID>IN_1</ID>1275 </input>
<output>
<ID>OUT</ID>1277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1573</ID>
<type>AA_AND2</type>
<position>145,250.5</position>
<input>
<ID>IN_0</ID>1276 </input>
<input>
<ID>IN_1</ID>1273 </input>
<output>
<ID>OUT</ID>1278 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1574</ID>
<type>AA_AND2</type>
<position>190.5,269</position>
<input>
<ID>IN_0</ID>1277 </input>
<input>
<ID>IN_1</ID>1279 </input>
<output>
<ID>OUT</ID>1281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1575</ID>
<type>AA_AND2</type>
<position>191,251.5</position>
<input>
<ID>IN_0</ID>1280 </input>
<input>
<ID>IN_1</ID>1278 </input>
<output>
<ID>OUT</ID>1282 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1576</ID>
<type>AE_DFF_LOW</type>
<position>149,217.5</position>
<input>
<ID>IN_0</ID>1275 </input>
<output>
<ID>OUT_0</ID>1287 </output>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1577</ID>
<type>AE_OR2</type>
<position>60.5,261</position>
<input>
<ID>IN_0</ID>1264 </input>
<input>
<ID>IN_1</ID>1265 </input>
<output>
<ID>OUT</ID>1302 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1578</ID>
<type>AE_DFF_LOW</type>
<position>195,217.5</position>
<input>
<ID>IN_0</ID>1279 </input>
<output>
<ID>OUT_0</ID>1288 </output>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1579</ID>
<type>AE_OR2</type>
<position>97,262</position>
<input>
<ID>IN_0</ID>1268 </input>
<input>
<ID>IN_1</ID>1270 </input>
<output>
<ID>OUT</ID>1305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1580</ID>
<type>AE_OR2</type>
<position>125.5,261.5</position>
<input>
<ID>IN_0</ID>1272 </input>
<input>
<ID>IN_1</ID>1273 </input>
<output>
<ID>OUT</ID>1306 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1581</ID>
<type>AE_OR2</type>
<position>154.5,261</position>
<input>
<ID>IN_0</ID>1277 </input>
<input>
<ID>IN_1</ID>1278 </input>
<output>
<ID>OUT</ID>1308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1582</ID>
<type>AE_OR2</type>
<position>198.5,260.5</position>
<input>
<ID>IN_0</ID>1281 </input>
<input>
<ID>IN_1</ID>1282 </input>
<output>
<ID>OUT</ID>1310 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1583</ID>
<type>AE_DFF_LOW</type>
<position>243,217</position>
<input>
<ID>IN_0</ID>1284 </input>
<output>
<ID>OUT_0</ID>1289 </output>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1584</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>247,237.5</position>
<input>
<ID>IN_0</ID>1262 </input>
<input>
<ID>IN_1</ID>1266 </input>
<input>
<ID>IN_2</ID>1271 </input>
<input>
<ID>IN_3</ID>1275 </input>
<input>
<ID>IN_4</ID>1279 </input>
<input>
<ID>IN_5</ID>1284 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1585</ID>
<type>AE_DFF_LOW</type>
<position>-33.5,253</position>
<input>
<ID>IN_0</ID>1317 </input>
<output>
<ID>OUTINV_0</ID>1319 </output>
<output>
<ID>OUT_0</ID>1318 </output>
<input>
<ID>clear</ID>1260 </input>
<input>
<ID>clock</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1587</ID>
<type>AE_OR2</type>
<position>542,35.5</position>
<input>
<ID>IN_0</ID>1387 </input>
<input>
<ID>IN_1</ID>1229 </input>
<output>
<ID>OUT</ID>1398 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1589</ID>
<type>AI_XOR2</type>
<position>526,33.5</position>
<input>
<ID>IN_0</ID>1249 </input>
<input>
<ID>IN_1</ID>1248 </input>
<output>
<ID>OUT</ID>1387 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1591</ID>
<type>GA_LED</type>
<position>563,35.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1595</ID>
<type>BA_NAND2</type>
<position>574,40.5</position>
<input>
<ID>IN_0</ID>1393 </input>
<input>
<ID>IN_1</ID>1399 </input>
<output>
<ID>OUT</ID>1397 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1601</ID>
<type>AO_XNOR2</type>
<position>554.5,33</position>
<input>
<ID>IN_0</ID>1398 </input>
<input>
<ID>IN_1</ID>1393 </input>
<output>
<ID>OUT</ID>1399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1409</ID>
<type>CC_PULSE</type>
<position>-81,258.5</position>
<output>
<ID>OUT_0</ID>1315 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1410</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>266.5,207</position>
<input>
<ID>IN_0</ID>1267 </input>
<input>
<ID>IN_1</ID>1285 </input>
<input>
<ID>IN_2</ID>1286 </input>
<input>
<ID>IN_3</ID>1287 </input>
<input>
<ID>IN_4</ID>1288 </input>
<input>
<ID>IN_5</ID>1289 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 10</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1411</ID>
<type>CC_PULSE</type>
<position>-79.5,240.5</position>
<output>
<ID>OUT_0</ID>1314 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1412</ID>
<type>EE_VDD</type>
<position>-29,293.5</position>
<output>
<ID>OUT_0</ID>1313 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1413</ID>
<type>AE_OR2</type>
<position>-42.5,241.5</position>
<input>
<ID>IN_0</ID>1315 </input>
<input>
<ID>IN_1</ID>1314 </input>
<output>
<ID>OUT</ID>1283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1414</ID>
<type>AE_DFF_LOW</type>
<position>465.5,61</position>
<input>
<ID>IN_0</ID>1231 </input>
<output>
<ID>OUT_0</ID>1237 </output>
<input>
<ID>clock</ID>1320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1415</ID>
<type>AE_SMALL_INVERTER</type>
<position>-60,258</position>
<input>
<ID>IN_0</ID>1315 </input>
<output>
<ID>OUT_0</ID>1316 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1609</ID>
<type>AA_TOGGLE</type>
<position>251.5,396</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1416</ID>
<type>AA_AND2</type>
<position>64,166.5</position>
<input>
<ID>IN_0</ID>1294 </input>
<input>
<ID>IN_1</ID>1293 </input>
<output>
<ID>OUT</ID>1295 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1417</ID>
<type>AI_XOR2</type>
<position>-45.5,254</position>
<input>
<ID>IN_0</ID>1314 </input>
<input>
<ID>IN_1</ID>1316 </input>
<output>
<ID>OUT</ID>1317 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1418</ID>
<type>AA_LABEL</type>
<position>-75.5,264.5</position>
<gparam>LABEL_TEXT Increment</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1419</ID>
<type>AA_AND2</type>
<position>138,180</position>
<input>
<ID>IN_0</ID>1296 </input>
<input>
<ID>IN_1</ID>1297 </input>
<output>
<ID>OUT</ID>1298 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1420</ID>
<type>AA_LABEL</type>
<position>-76.5,235.5</position>
<gparam>LABEL_TEXT Decrement</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1421</ID>
<type>AA_AND2</type>
<position>201,181.5</position>
<input>
<ID>IN_0</ID>1299 </input>
<input>
<ID>IN_1</ID>1300 </input>
<output>
<ID>OUT</ID>1301 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1422</ID>
<type>AI_XOR2</type>
<position>14.5,272.5</position>
<input>
<ID>IN_0</ID>1290 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1292 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1423</ID>
<type>AE_DFF_LOW</type>
<position>479,61</position>
<input>
<ID>IN_0</ID>1232 </input>
<output>
<ID>OUT_0</ID>1238 </output>
<input>
<ID>clock</ID>1320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1424</ID>
<type>AI_XOR2</type>
<position>65.5,275</position>
<input>
<ID>IN_0</ID>1302 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1303 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1425</ID>
<type>AI_XOR2</type>
<position>102,275.5</position>
<input>
<ID>IN_0</ID>1305 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1304 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1426</ID>
<type>AI_XOR2</type>
<position>130.5,275</position>
<input>
<ID>IN_0</ID>1306 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1307 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1427</ID>
<type>AI_XOR2</type>
<position>160.5,275</position>
<input>
<ID>IN_0</ID>1308 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1309 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1428</ID>
<type>AI_XOR2</type>
<position>208,277</position>
<input>
<ID>IN_0</ID>1310 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1311 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1429</ID>
<type>AA_AND4</type>
<position>42.5,144.5</position>
<input>
<ID>IN_0</ID>1301 </input>
<input>
<ID>IN_1</ID>1298 </input>
<input>
<ID>IN_2</ID>1295 </input>
<input>
<ID>IN_3</ID>1319 </input>
<output>
<ID>OUT</ID>1291 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1430</ID>
<type>AE_DFF_LOW</type>
<position>494,61</position>
<input>
<ID>IN_0</ID>1233 </input>
<output>
<ID>OUT_0</ID>1239 </output>
<input>
<ID>clock</ID>1320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1431</ID>
<type>AA_INVERTER</type>
<position>58,189.5</position>
<input>
<ID>IN_0</ID>1262 </input>
<output>
<ID>OUT_0</ID>1293 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1432</ID>
<type>AA_INVERTER</type>
<position>70.5,188.5</position>
<input>
<ID>IN_0</ID>1266 </input>
<output>
<ID>OUT_0</ID>1294 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1433</ID>
<type>AA_INVERTER</type>
<position>134.5,189.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<output>
<ID>OUT_0</ID>1297 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1434</ID>
<type>AA_INVERTER</type>
<position>141.5,189.5</position>
<input>
<ID>IN_0</ID>1275 </input>
<output>
<ID>OUT_0</ID>1296 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1435</ID>
<type>AE_DFF_LOW</type>
<position>504.5,61</position>
<input>
<ID>IN_0</ID>1234 </input>
<output>
<ID>OUT_0</ID>1240 </output>
<input>
<ID>clock</ID>1320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1436</ID>
<type>AA_INVERTER</type>
<position>199,190</position>
<input>
<ID>IN_0</ID>1279 </input>
<output>
<ID>OUT_0</ID>1300 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1437</ID>
<type>AA_INVERTER</type>
<position>204.5,190.5</position>
<input>
<ID>IN_0</ID>1284 </input>
<output>
<ID>OUT_0</ID>1299 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1438</ID>
<type>AA_LABEL</type>
<position>266.5,197</position>
<gparam>LABEL_TEXT Actual Timer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1439</ID>
<type>AA_AND2</type>
<position>-36,287</position>
<input>
<ID>IN_0</ID>1313 </input>
<input>
<ID>IN_1</ID>1312 </input>
<output>
<ID>OUT</ID>1290 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1440</ID>
<type>AA_LABEL</type>
<position>93,296.5</position>
<gparam>LABEL_TEXT Setting Mode</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1441</ID>
<type>AE_DFF_LOW</type>
<position>517.5,61</position>
<input>
<ID>IN_0</ID>1235 </input>
<output>
<ID>OUT_0</ID>1241 </output>
<input>
<ID>clock</ID>1320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1442</ID>
<type>AA_LABEL</type>
<position>-42,300</position>
<gparam>LABEL_TEXT On/Off- Settings/Cycle</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1444</ID>
<type>AA_LABEL</type>
<position>-55.5,488.5</position>
<gparam>LABEL_TEXT Water Button</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1445</ID>
<type>AE_SMALL_INVERTER</type>
<position>456.5,53.5</position>
<input>
<ID>IN_0</ID>1236 </input>
<output>
<ID>OUT_0</ID>1242 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1446</ID>
<type>AA_LABEL</type>
<position>95,447.5</position>
<gparam>LABEL_TEXT Buffer Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1447</ID>
<type>AA_LABEL</type>
<position>37,499</position>
<gparam>LABEL_TEXT Seconds Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1448</ID>
<type>AE_SMALL_INVERTER</type>
<position>471.5,53.5</position>
<input>
<ID>IN_0</ID>1237 </input>
<output>
<ID>OUT_0</ID>1243 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1449</ID>
<type>BE_JKFF_LOW_NT</type>
<position>224,386</position>
<input>
<ID>J</ID>1370 </input>
<input>
<ID>K</ID>1390 </input>
<output>
<ID>Q</ID>1407 </output>
<input>
<ID>clear</ID>1397 </input>
<input>
<ID>clock</ID>1320 </input>
<output>
<ID>nQ</ID>1408 </output>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1450</ID>
<type>AA_LABEL</type>
<position>93.5,426</position>
<gparam>LABEL_TEXT Actual Seconds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1451</ID>
<type>AE_SMALL_INVERTER</type>
<position>486.5,53.5</position>
<input>
<ID>IN_0</ID>1238 </input>
<output>
<ID>OUT_0</ID>1244 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1452</ID>
<type>AA_LABEL</type>
<position>167.5,407.5</position>
<gparam>LABEL_TEXT Minutes Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1453</ID>
<type>AE_SMALL_INVERTER</type>
<position>498,54</position>
<input>
<ID>IN_0</ID>1239 </input>
<output>
<ID>OUT_0</ID>1245 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1454</ID>
<type>AA_LABEL</type>
<position>230.5,372</position>
<gparam>LABEL_TEXT Buffer Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1455</ID>
<type>AE_SMALL_INVERTER</type>
<position>511,53.5</position>
<input>
<ID>IN_0</ID>1240 </input>
<output>
<ID>OUT_0</ID>1246 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1456</ID>
<type>AI_XOR2</type>
<position>109.5,472</position>
<input>
<ID>IN_0</ID>1408 </input>
<input>
<ID>IN_1</ID>1329 </input>
<output>
<ID>OUT</ID>1335 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1457</ID>
<type>AA_LABEL</type>
<position>114,482</position>
<gparam>LABEL_TEXT Both on seconds counter stop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1458</ID>
<type>AE_SMALL_INVERTER</type>
<position>524,54</position>
<input>
<ID>IN_0</ID>1241 </input>
<output>
<ID>OUT_0</ID>1247 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1459</ID>
<type>AA_LABEL</type>
<position>240,343</position>
<gparam>LABEL_TEXT Actual Minutes</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1460</ID>
<type>AI_XOR2</type>
<position>208.5,384</position>
<input>
<ID>IN_0</ID>1336 </input>
<input>
<ID>IN_1</ID>1407 </input>
<output>
<ID>OUT</ID>1324 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1461</ID>
<type>AA_INVERTER</type>
<position>217.5,401</position>
<input>
<ID>IN_0</ID>1330 </input>
<output>
<ID>OUT_0</ID>1390 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1462</ID>
<type>AA_AND2</type>
<position>-29,448.5</position>
<input>
<ID>IN_0</ID>1370 </input>
<input>
<ID>IN_1</ID>1320 </input>
<output>
<ID>OUT</ID>1342 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1463</ID>
<type>AA_LABEL</type>
<position>-40,374.5</position>
<gparam>LABEL_TEXT Abort</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1464</ID>
<type>AE_OR2</type>
<position>24.5,392.5</position>
<input>
<ID>IN_0</ID>1353 </input>
<input>
<ID>IN_1</ID>1352 </input>
<output>
<ID>OUT</ID>1325 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1465</ID>
<type>AA_TOGGLE</type>
<position>-38,379.5</position>
<output>
<ID>OUT_0</ID>1336 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1466</ID>
<type>AE_OR4</type>
<position>-7.5,401</position>
<input>
<ID>IN_0</ID>1351 </input>
<input>
<ID>IN_1</ID>1350 </input>
<input>
<ID>IN_2</ID>1349 </input>
<input>
<ID>IN_3</ID>1348 </input>
<output>
<ID>OUT</ID>1322 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1467</ID>
<type>AE_OR2</type>
<position>-21.5,395.5</position>
<input>
<ID>IN_0</ID>1325 </input>
<input>
<ID>IN_1</ID>1322 </input>
<output>
<ID>OUT</ID>1332 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1468</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-16.5,461</position>
<input>
<ID>J</ID>1370 </input>
<input>
<ID>K</ID>1370 </input>
<output>
<ID>Q</ID>1341 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1469</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-3,461</position>
<input>
<ID>J</ID>1341 </input>
<input>
<ID>K</ID>1341 </input>
<output>
<ID>Q</ID>1343 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1470</ID>
<type>AA_AND2</type>
<position>-28,405</position>
<input>
<ID>IN_0</ID>1324 </input>
<input>
<ID>IN_1</ID>1370 </input>
<output>
<ID>OUT</ID>1326 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1471</ID>
<type>BE_JKFF_LOW_NT</type>
<position>13,461</position>
<input>
<ID>J</ID>1337 </input>
<input>
<ID>K</ID>1337 </input>
<output>
<ID>Q</ID>1345 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1472</ID>
<type>AA_TOGGLE</type>
<position>326,169.5</position>
<output>
<ID>OUT_0</ID>1229 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1473</ID>
<type>AE_OR2</type>
<position>-46.5,408</position>
<input>
<ID>IN_0</ID>1333 </input>
<input>
<ID>IN_1</ID>1326 </input>
<output>
<ID>OUT</ID>1334 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1474</ID>
<type>BE_JKFF_LOW_NT</type>
<position>29,460.5</position>
<input>
<ID>J</ID>1338 </input>
<input>
<ID>K</ID>1338 </input>
<output>
<ID>Q</ID>1344 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1475</ID>
<type>AA_AND4</type>
<position>474.5,37</position>
<input>
<ID>IN_0</ID>1245 </input>
<input>
<ID>IN_1</ID>1244 </input>
<input>
<ID>IN_2</ID>1243 </input>
<input>
<ID>IN_3</ID>1242 </input>
<output>
<ID>OUT</ID>1248 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1476</ID>
<type>BE_JKFF_LOW_NT</type>
<position>45,460</position>
<input>
<ID>J</ID>1339 </input>
<input>
<ID>K</ID>1339 </input>
<output>
<ID>Q</ID>1346 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1477</ID>
<type>BE_JKFF_LOW_NT</type>
<position>62,460</position>
<input>
<ID>J</ID>1340 </input>
<input>
<ID>K</ID>1340 </input>
<output>
<ID>Q</ID>1347 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1478</ID>
<type>AI_XOR2</type>
<position>94.5,463</position>
<input>
<ID>IN_0</ID>1336 </input>
<input>
<ID>IN_1</ID>1335 </input>
<output>
<ID>OUT</ID>1328 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1479</ID>
<type>AA_TOGGLE</type>
<position>-44,481.5</position>
<output>
<ID>OUT_0</ID>1409 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1480</ID>
<type>AA_LABEL</type>
<position>-60,415</position>
<gparam>LABEL_TEXT Water On/Off</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1481</ID>
<type>BE_JKFF_LOW_NT</type>
<position>112,388</position>
<input>
<ID>J</ID>1370 </input>
<input>
<ID>K</ID>1370 </input>
<output>
<ID>Q</ID>1358 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1482</ID>
<type>AA_AND2</type>
<position>-39,396.5</position>
<input>
<ID>IN_0</ID>1332 </input>
<input>
<ID>IN_1</ID>1370 </input>
<output>
<ID>OUT</ID>1333 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1483</ID>
<type>BE_JKFF_LOW_NT</type>
<position>125.5,388</position>
<input>
<ID>J</ID>1358 </input>
<input>
<ID>K</ID>1358 </input>
<output>
<ID>Q</ID>1359 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1484</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>79.5,446.5</position>
<input>
<ID>IN_0</ID>1341 </input>
<input>
<ID>IN_1</ID>1343 </input>
<input>
<ID>IN_2</ID>1345 </input>
<input>
<ID>IN_3</ID>1344 </input>
<input>
<ID>IN_4</ID>1346 </input>
<input>
<ID>IN_5</ID>1347 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1485</ID>
<type>BE_JKFF_LOW_NT</type>
<position>141.5,388</position>
<input>
<ID>J</ID>1354 </input>
<input>
<ID>K</ID>1354 </input>
<output>
<ID>Q</ID>1361 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1486</ID>
<type>AA_AND2</type>
<position>511,38</position>
<input>
<ID>IN_0</ID>1247 </input>
<input>
<ID>IN_1</ID>1246 </input>
<output>
<ID>OUT</ID>1249 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1487</ID>
<type>GA_LED</type>
<position>-58.5,408</position>
<input>
<ID>N_in1</ID>1334 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1488</ID>
<type>BE_JKFF_LOW_NT</type>
<position>157.5,387.5</position>
<input>
<ID>J</ID>1355 </input>
<input>
<ID>K</ID>1355 </input>
<output>
<ID>Q</ID>1360 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1489</ID>
<type>AA_AND2</type>
<position>490,25</position>
<input>
<ID>IN_0</ID>1249 </input>
<input>
<ID>IN_1</ID>1248 </input>
<output>
<ID>OUT</ID>1393 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1490</ID>
<type>AA_LABEL</type>
<position>-8,390</position>
<gparam>LABEL_TEXT Output of Flip-flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1491</ID>
<type>BE_JKFF_LOW_NT</type>
<position>173.5,388</position>
<input>
<ID>J</ID>1356 </input>
<input>
<ID>K</ID>1356 </input>
<output>
<ID>Q</ID>1362 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1492</ID>
<type>BB_CLOCK</type>
<position>-43.5,447.5</position>
<output>
<ID>CLK</ID>1320 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 3</lparam></gate>
<gate>
<ID>1493</ID>
<type>BE_JKFF_LOW_NT</type>
<position>190.5,388</position>
<input>
<ID>J</ID>1357 </input>
<input>
<ID>K</ID>1357 </input>
<output>
<ID>Q</ID>1363 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1494</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>202.5,373.5</position>
<input>
<ID>IN_0</ID>1358 </input>
<input>
<ID>IN_1</ID>1359 </input>
<input>
<ID>IN_2</ID>1361 </input>
<input>
<ID>IN_3</ID>1360 </input>
<input>
<ID>IN_4</ID>1362 </input>
<input>
<ID>IN_5</ID>1363 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1495</ID>
<type>AA_AND2</type>
<position>4,471.5</position>
<input>
<ID>IN_0</ID>1341 </input>
<input>
<ID>IN_1</ID>1343 </input>
<output>
<ID>OUT</ID>1337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1496</ID>
<type>AI_XOR2</type>
<position>-34.5,473.5</position>
<input>
<ID>IN_0</ID>1397 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1497</ID>
<type>AA_AND2</type>
<position>132.5,398.5</position>
<input>
<ID>IN_0</ID>1358 </input>
<input>
<ID>IN_1</ID>1359 </input>
<output>
<ID>OUT</ID>1354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1498</ID>
<type>AA_AND2</type>
<position>149.5,397.5</position>
<input>
<ID>IN_0</ID>1354 </input>
<input>
<ID>IN_1</ID>1361 </input>
<output>
<ID>OUT</ID>1355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1499</ID>
<type>AA_AND2</type>
<position>21,470.5</position>
<input>
<ID>IN_0</ID>1337 </input>
<input>
<ID>IN_1</ID>1345 </input>
<output>
<ID>OUT</ID>1338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1500</ID>
<type>AA_AND2</type>
<position>164.5,396.5</position>
<input>
<ID>IN_0</ID>1355 </input>
<input>
<ID>IN_1</ID>1360 </input>
<output>
<ID>OUT</ID>1356 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1501</ID>
<type>AA_AND2</type>
<position>182,395.5</position>
<input>
<ID>IN_0</ID>1356 </input>
<input>
<ID>IN_1</ID>1362 </input>
<output>
<ID>OUT</ID>1357 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1502</ID>
<type>AA_AND2</type>
<position>36,469.5</position>
<input>
<ID>IN_0</ID>1338 </input>
<input>
<ID>IN_1</ID>1344 </input>
<output>
<ID>OUT</ID>1339 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1503</ID>
<type>BA_NAND4</type>
<position>204,398.5</position>
<input>
<ID>IN_0</ID>1361 </input>
<input>
<ID>IN_1</ID>1360 </input>
<input>
<ID>IN_2</ID>1362 </input>
<input>
<ID>IN_3</ID>1363 </input>
<output>
<ID>OUT</ID>1330 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1504</ID>
<type>AE_DFF_LOW</type>
<position>121,353</position>
<input>
<ID>IN_0</ID>1358 </input>
<output>
<ID>OUT_0</ID>1364 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1505</ID>
<type>AA_AND2</type>
<position>53.5,468.5</position>
<input>
<ID>IN_0</ID>1339 </input>
<input>
<ID>IN_1</ID>1346 </input>
<output>
<ID>OUT</ID>1340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1506</ID>
<type>AE_DFF_LOW</type>
<position>137.5,353</position>
<input>
<ID>IN_0</ID>1359 </input>
<output>
<ID>OUT_0</ID>1365 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1507</ID>
<type>AE_DFF_LOW</type>
<position>152,353</position>
<input>
<ID>IN_0</ID>1361 </input>
<output>
<ID>OUT_0</ID>1366 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1508</ID>
<type>BA_NAND4</type>
<position>75.5,471.5</position>
<input>
<ID>IN_0</ID>1345 </input>
<input>
<ID>IN_1</ID>1344 </input>
<input>
<ID>IN_2</ID>1346 </input>
<input>
<ID>IN_3</ID>1347 </input>
<output>
<ID>OUT</ID>1329 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1509</ID>
<type>AE_DFF_LOW</type>
<position>169,353</position>
<input>
<ID>IN_0</ID>1360 </input>
<output>
<ID>OUT_0</ID>1367 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1510</ID>
<type>AE_DFF_LOW</type>
<position>185,353</position>
<input>
<ID>IN_0</ID>1362 </input>
<output>
<ID>OUT_0</ID>1368 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1511</ID>
<type>AE_DFF_LOW</type>
<position>203,353</position>
<input>
<ID>IN_0</ID>1363 </input>
<output>
<ID>OUT_0</ID>1369 </output>
<input>
<ID>clear</ID>1324 </input>
<input>
<ID>clock</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1512</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>223,343.5</position>
<input>
<ID>IN_0</ID>1364 </input>
<input>
<ID>IN_1</ID>1365 </input>
<input>
<ID>IN_2</ID>1366 </input>
<input>
<ID>IN_3</ID>1367 </input>
<input>
<ID>IN_4</ID>1368 </input>
<input>
<ID>IN_5</ID>1369 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1513</ID>
<type>AA_INVERTER</type>
<position>110.5,446</position>
<input>
<ID>IN_0</ID>1328 </input>
<output>
<ID>OUT_0</ID>1371 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1514</ID>
<type>AE_DFF_LOW</type>
<position>-7.5,426</position>
<input>
<ID>IN_0</ID>1341 </input>
<output>
<ID>OUT_0</ID>1348 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1515</ID>
<type>AE_DFF_LOW</type>
<position>9,426</position>
<input>
<ID>IN_0</ID>1343 </input>
<output>
<ID>OUT_0</ID>1349 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1516</ID>
<type>AE_DFF_LOW</type>
<position>23.5,426</position>
<input>
<ID>IN_0</ID>1345 </input>
<output>
<ID>OUT_0</ID>1350 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1517</ID>
<type>AE_DFF_LOW</type>
<position>40.5,426</position>
<input>
<ID>IN_0</ID>1344 </input>
<output>
<ID>OUT_0</ID>1351 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1518</ID>
<type>AE_DFF_LOW</type>
<position>56.5,426</position>
<input>
<ID>IN_0</ID>1346 </input>
<output>
<ID>OUT_0</ID>1352 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1519</ID>
<type>AE_DFF_LOW</type>
<position>74.5,426</position>
<input>
<ID>IN_0</ID>1347 </input>
<output>
<ID>OUT_0</ID>1353 </output>
<input>
<ID>clear</ID>1328 </input>
<input>
<ID>clock</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1520</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>94.5,416.5</position>
<input>
<ID>IN_0</ID>1348 </input>
<input>
<ID>IN_1</ID>1349 </input>
<input>
<ID>IN_2</ID>1350 </input>
<input>
<ID>IN_3</ID>1351 </input>
<input>
<ID>IN_4</ID>1352 </input>
<input>
<ID>IN_5</ID>1353 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1521</ID>
<type>AA_AND2</type>
<position>-43,457</position>
<input>
<ID>IN_0</ID>1409 </input>
<input>
<ID>IN_1</ID>1258 </input>
<output>
<ID>OUT</ID>1370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1522</ID>
<type>AE_DFF_LOW</type>
<position>-99,290</position>
<input>
<ID>IN_0</ID>1253 </input>
<output>
<ID>OUTINV_0</ID>1259 </output>
<output>
<ID>OUT_0</ID>1257 </output>
<input>
<ID>clock</ID>1255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1523</ID>
<type>AA_TOGGLE</type>
<position>-111.5,292</position>
<output>
<ID>OUT_0</ID>1253 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1524</ID>
<type>AI_XOR2</type>
<position>445.5,70</position>
<input>
<ID>IN_0</ID>1364 </input>
<input>
<ID>IN_1</ID>1373 </input>
<output>
<ID>OUT</ID>1230 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1525</ID>
<type>AI_XOR2</type>
<position>459,70</position>
<input>
<ID>IN_0</ID>1365 </input>
<input>
<ID>IN_1</ID>1375 </input>
<output>
<ID>OUT</ID>1231 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1526</ID>
<type>AA_AND2</type>
<position>-82.5,301</position>
<input>
<ID>IN_0</ID>1257 </input>
<input>
<ID>IN_1</ID>1256 </input>
<output>
<ID>OUT</ID>1258 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1527</ID>
<type>AI_XOR2</type>
<position>472,70</position>
<input>
<ID>IN_0</ID>1366 </input>
<input>
<ID>IN_1</ID>1377 </input>
<output>
<ID>OUT</ID>1232 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1528</ID>
<type>AI_XOR2</type>
<position>485,70</position>
<input>
<ID>IN_0</ID>1367 </input>
<input>
<ID>IN_1</ID>1379 </input>
<output>
<ID>OUT</ID>1233 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1529</ID>
<type>AI_XOR2</type>
<position>497.5,69.5</position>
<input>
<ID>IN_0</ID>1368 </input>
<input>
<ID>IN_1</ID>1381 </input>
<output>
<ID>OUT</ID>1234 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1530</ID>
<type>AE_SMALL_INVERTER</type>
<position>-88.5,289</position>
<input>
<ID>IN_0</ID>1259 </input>
<output>
<ID>OUT_0</ID>1260 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1531</ID>
<type>AI_XOR2</type>
<position>510,69.5</position>
<input>
<ID>IN_0</ID>1369 </input>
<input>
<ID>IN_1</ID>1383 </input>
<output>
<ID>OUT</ID>1235 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1532</ID>
<type>AA_LABEL</type>
<position>39.5,279.5</position>
<gparam>LABEL_TEXT Default Power</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1533</ID>
<type>AE_DFF_LOW</type>
<position>-49,288</position>
<input>
<ID>IN_0</ID>1254 </input>
<output>
<ID>OUTINV_0</ID>1256 </output>
<output>
<ID>OUT_0</ID>1312 </output>
<input>
<ID>clear</ID>1260 </input>
<input>
<ID>clock</ID>1255 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1534</ID>
<type>BB_CLOCK</type>
<position>-64,284.5</position>
<output>
<ID>CLK</ID>1255 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1535</ID>
<type>AA_TOGGLE</type>
<position>332,23.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1536</ID>
<type>AA_LABEL</type>
<position>337,173</position>
<gparam>LABEL_TEXT Zone 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1537</ID>
<type>AA_LABEL</type>
<position>337,18</position>
<gparam>LABEL_TEXT Zone 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1538</ID>
<type>BE_JKFF_LOW_NT</type>
<position>424.5,107</position>
<input>
<ID>J</ID>1372 </input>
<output>
<ID>Q</ID>1373 </output>
<input>
<ID>clear</ID>1385 </input>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1539</ID>
<type>BE_JKFF_LOW_NT</type>
<position>411.5,117</position>
<input>
<ID>J</ID>1374 </input>
<output>
<ID>Q</ID>1375 </output>
<input>
<ID>clear</ID>1385 </input>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1540</ID>
<type>BE_JKFF_LOW_NT</type>
<position>398.5,128</position>
<input>
<ID>J</ID>1376 </input>
<output>
<ID>Q</ID>1377 </output>
<input>
<ID>clear</ID>1385 </input>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1541</ID>
<type>BE_JKFF_LOW_NT</type>
<position>391,137</position>
<input>
<ID>J</ID>1378 </input>
<output>
<ID>Q</ID>1379 </output>
<input>
<ID>clear</ID>1385 </input>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1542</ID>
<type>BE_JKFF_LOW_NT</type>
<position>382.5,144.5</position>
<input>
<ID>J</ID>1380 </input>
<output>
<ID>Q</ID>1381 </output>
<input>
<ID>clear</ID>1385 </input>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1543</ID>
<type>BE_JKFF_LOW_NT</type>
<position>373.5,152</position>
<input>
<ID>J</ID>1382 </input>
<output>
<ID>Q</ID>1383 </output>
<input>
<ID>clear</ID>1385 </input>
<input>
<ID>clock</ID>1384 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>1351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,416.5,89.5,416.5</points>
<connection>
<GID>1520</GID>
<name>IN_3</name></connection>
<intersection>46 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46,398,46,428</points>
<intersection>398 8</intersection>
<intersection>416.5 1</intersection>
<intersection>428 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,428,46,428</points>
<connection>
<GID>1517</GID>
<name>OUT_0</name></connection>
<intersection>46 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-4.5,398,46,398</points>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection>
<intersection>46 3</intersection></hsegment></shape></wire>
<wire>
<ID>1352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,417.5,89.5,417.5</points>
<connection>
<GID>1520</GID>
<name>IN_4</name></connection>
<intersection>27.5 7</intersection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,417.5,60.5,428</points>
<intersection>417.5 1</intersection>
<intersection>428 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>59.5,428,60.5,428</points>
<connection>
<GID>1518</GID>
<name>OUT_0</name></connection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>27.5,393.5,27.5,417.5</points>
<connection>
<GID>1464</GID>
<name>IN_1</name></connection>
<intersection>417.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80.5,418.5,89.5,418.5</points>
<connection>
<GID>1520</GID>
<name>IN_5</name></connection>
<intersection>80.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>80.5,391.5,80.5,428</points>
<intersection>391.5 8</intersection>
<intersection>418.5 1</intersection>
<intersection>428 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>77.5,428,80.5,428</points>
<connection>
<GID>1519</GID>
<name>OUT_0</name></connection>
<intersection>80.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>27.5,391.5,80.5,391.5</points>
<connection>
<GID>1464</GID>
<name>IN_0</name></connection>
<intersection>80.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,386,137,398.5</points>
<intersection>386 4</intersection>
<intersection>390 2</intersection>
<intersection>398.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,398.5,146.5,398.5</points>
<connection>
<GID>1497</GID>
<name>OUT</name></connection>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137,390,138.5,390</points>
<connection>
<GID>1485</GID>
<name>J</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>137,386,138.5,386</points>
<connection>
<GID>1485</GID>
<name>K</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>1355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,385.5,153.5,397.5</points>
<intersection>385.5 4</intersection>
<intersection>389.5 2</intersection>
<intersection>397.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,397.5,161.5,397.5</points>
<connection>
<GID>1498</GID>
<name>OUT</name></connection>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<intersection>153.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153.5,389.5,154.5,389.5</points>
<connection>
<GID>1488</GID>
<name>J</name></connection>
<intersection>153.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>153.5,385.5,154.5,385.5</points>
<connection>
<GID>1488</GID>
<name>K</name></connection>
<intersection>153.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,386,169,396.5</points>
<intersection>386 4</intersection>
<intersection>390 2</intersection>
<intersection>396.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,396.5,179,396.5</points>
<connection>
<GID>1500</GID>
<name>OUT</name></connection>
<connection>
<GID>1501</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,390,170.5,390</points>
<connection>
<GID>1491</GID>
<name>J</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>169,386,170.5,386</points>
<connection>
<GID>1491</GID>
<name>K</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>1357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,386,186,395.5</points>
<intersection>386 4</intersection>
<intersection>390 2</intersection>
<intersection>395.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,395.5,186,395.5</points>
<connection>
<GID>1501</GID>
<name>OUT</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,390,187.5,390</points>
<connection>
<GID>1493</GID>
<name>J</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>186,386,187.5,386</points>
<connection>
<GID>1493</GID>
<name>K</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire>
<wire>
<ID>1358</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,390,122.5,390</points>
<connection>
<GID>1481</GID>
<name>Q</name></connection>
<connection>
<GID>1483</GID>
<name>J</name></connection>
<intersection>116 3</intersection>
<intersection>118.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,355,116,390</points>
<intersection>355 10</intersection>
<intersection>370.5 4</intersection>
<intersection>386 9</intersection>
<intersection>390 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>116,370.5,197.5,370.5</points>
<connection>
<GID>1494</GID>
<name>IN_0</name></connection>
<intersection>116 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>118.5,390,118.5,399.5</points>
<intersection>390 1</intersection>
<intersection>399.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>118.5,399.5,129.5,399.5</points>
<connection>
<GID>1497</GID>
<name>IN_0</name></connection>
<intersection>118.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116,386,122.5,386</points>
<connection>
<GID>1483</GID>
<name>K</name></connection>
<intersection>116 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116,355,118,355</points>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>116 3</intersection></hsegment></shape></wire>
<wire>
<ID>1359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,355,129.5,397.5</points>
<connection>
<GID>1497</GID>
<name>IN_1</name></connection>
<intersection>355 8</intersection>
<intersection>371.5 1</intersection>
<intersection>390 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,371.5,197.5,371.5</points>
<connection>
<GID>1494</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>128.5,390,129.5,390</points>
<connection>
<GID>1483</GID>
<name>Q</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>129.5,355,134.5,355</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,373.5,197.5,373.5</points>
<connection>
<GID>1494</GID>
<name>IN_3</name></connection>
<intersection>161.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>161.5,355,161.5,399.5</points>
<connection>
<GID>1500</GID>
<name>IN_1</name></connection>
<intersection>355 9</intersection>
<intersection>373.5 1</intersection>
<intersection>389.5 4</intersection>
<intersection>399.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>160.5,389.5,161.5,389.5</points>
<connection>
<GID>1488</GID>
<name>Q</name></connection>
<intersection>161.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>161.5,399.5,201,399.5</points>
<connection>
<GID>1503</GID>
<name>IN_1</name></connection>
<intersection>161.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>161.5,355,166,355</points>
<connection>
<GID>1509</GID>
<name>IN_0</name></connection>
<intersection>161.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,355,145.5,401.5</points>
<intersection>355 9</intersection>
<intersection>372.5 4</intersection>
<intersection>390 3</intersection>
<intersection>396.5 2</intersection>
<intersection>401.5 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>145.5,396.5,146.5,396.5</points>
<connection>
<GID>1498</GID>
<name>IN_1</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>144.5,390,145.5,390</points>
<connection>
<GID>1485</GID>
<name>Q</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>145.5,372.5,197.5,372.5</points>
<connection>
<GID>1494</GID>
<name>IN_2</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>145.5,401.5,201,401.5</points>
<connection>
<GID>1503</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>145.5,355,149,355</points>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,355,177.5,397.5</points>
<intersection>355 8</intersection>
<intersection>374.5 3</intersection>
<intersection>390 1</intersection>
<intersection>397.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176.5,390,177.5,390</points>
<connection>
<GID>1491</GID>
<name>Q</name></connection>
<intersection>177.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177.5,397.5,201,397.5</points>
<connection>
<GID>1503</GID>
<name>IN_2</name></connection>
<intersection>177.5 0</intersection>
<intersection>179 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>177.5,374.5,197.5,374.5</points>
<connection>
<GID>1494</GID>
<name>IN_4</name></connection>
<intersection>177.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>179,394.5,179,397.5</points>
<connection>
<GID>1501</GID>
<name>IN_1</name></connection>
<intersection>397.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>177.5,355,182,355</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<intersection>177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,355,195.5,395.5</points>
<intersection>355 5</intersection>
<intersection>375.5 2</intersection>
<intersection>390 1</intersection>
<intersection>395.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,390,195.5,390</points>
<connection>
<GID>1493</GID>
<name>Q</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195.5,375.5,197.5,375.5</points>
<connection>
<GID>1494</GID>
<name>IN_5</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>195.5,395.5,201,395.5</points>
<connection>
<GID>1503</GID>
<name>IN_3</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>195.5,355,200,355</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125.5,303,439,303</points>
<intersection>125.5 3</intersection>
<intersection>439 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>125.5,303,125.5,355</points>
<intersection>303 1</intersection>
<intersection>340.5 7</intersection>
<intersection>355 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124,355,125.5,355</points>
<connection>
<GID>1504</GID>
<name>OUT_0</name></connection>
<intersection>125.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>439,76,439,303</points>
<intersection>76 11</intersection>
<intersection>303 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>125.5,340.5,218,340.5</points>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection>
<intersection>125.5 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>439,76,446.5,76</points>
<intersection>439 5</intersection>
<intersection>446.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>446.5,73,446.5,76</points>
<connection>
<GID>1524</GID>
<name>IN_0</name></connection>
<intersection>76 11</intersection></vsegment></shape></wire>
<wire>
<ID>1365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,307.5,460,307.5</points>
<intersection>142 3</intersection>
<intersection>460 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>142,307.5,142,355</points>
<intersection>307.5 1</intersection>
<intersection>341.5 7</intersection>
<intersection>355 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>140.5,355,142,355</points>
<connection>
<GID>1506</GID>
<name>OUT_0</name></connection>
<intersection>142 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>460,73,460,307.5</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<intersection>307.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>142,341.5,218,341.5</points>
<connection>
<GID>1512</GID>
<name>IN_1</name></connection>
<intersection>142 3</intersection></hsegment></shape></wire>
<wire>
<ID>1366</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,312,474,312</points>
<intersection>156 3</intersection>
<intersection>474 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>156,312,156,355</points>
<intersection>312 1</intersection>
<intersection>342.5 7</intersection>
<intersection>355 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>155,355,156,355</points>
<connection>
<GID>1507</GID>
<name>OUT_0</name></connection>
<intersection>156 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>474,73,474,312</points>
<intersection>73 9</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>156,342.5,218,342.5</points>
<connection>
<GID>1512</GID>
<name>IN_2</name></connection>
<intersection>156 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>473,73,474,73</points>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection>
<intersection>474 5</intersection></hsegment></shape></wire>
<wire>
<ID>1367</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174.5,316.5,487,316.5</points>
<intersection>174.5 3</intersection>
<intersection>487 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>174.5,316.5,174.5,355</points>
<intersection>316.5 1</intersection>
<intersection>343.5 7</intersection>
<intersection>355 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172,355,174.5,355</points>
<connection>
<GID>1509</GID>
<name>OUT_0</name></connection>
<intersection>174.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>487,73,487,316.5</points>
<intersection>73 9</intersection>
<intersection>316.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>174.5,343.5,218,343.5</points>
<connection>
<GID>1512</GID>
<name>IN_3</name></connection>
<intersection>174.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>486,73,487,73</points>
<connection>
<GID>1528</GID>
<name>IN_0</name></connection>
<intersection>487 5</intersection></hsegment></shape></wire>
<wire>
<ID>1368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,319.5,499.5,319.5</points>
<intersection>189.5 3</intersection>
<intersection>499.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>189.5,319.5,189.5,355</points>
<intersection>319.5 1</intersection>
<intersection>344.5 7</intersection>
<intersection>355 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>188,355,189.5,355</points>
<connection>
<GID>1510</GID>
<name>OUT_0</name></connection>
<intersection>189.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>499.5,72.5,499.5,319.5</points>
<intersection>72.5 9</intersection>
<intersection>319.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>189.5,344.5,218,344.5</points>
<connection>
<GID>1512</GID>
<name>IN_4</name></connection>
<intersection>189.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>498.5,72.5,499.5,72.5</points>
<connection>
<GID>1529</GID>
<name>IN_0</name></connection>
<intersection>499.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,324.5,212,355</points>
<intersection>324.5 5</intersection>
<intersection>345.5 8</intersection>
<intersection>355 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206,355,212,355</points>
<connection>
<GID>1511</GID>
<name>OUT_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>212,324.5,512,324.5</points>
<intersection>212 0</intersection>
<intersection>512 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>512,72.5,512,324.5</points>
<intersection>72.5 10</intersection>
<intersection>324.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>212,345.5,218,345.5</points>
<connection>
<GID>1512</GID>
<name>IN_5</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>511,72.5,512,72.5</points>
<connection>
<GID>1531</GID>
<name>IN_0</name></connection>
<intersection>512 6</intersection></hsegment></shape></wire>
<wire>
<ID>1370</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>105.5,386,105.5,415</points>
<intersection>386 4</intersection>
<intersection>390 17</intersection>
<intersection>415 31</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-33.5,386,109,386</points>
<connection>
<GID>1481</GID>
<name>K</name></connection>
<intersection>-33.5 11</intersection>
<intersection>105.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-33.5,463,-19.5,463</points>
<connection>
<GID>1468</GID>
<name>J</name></connection>
<intersection>-33.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-33.5,386,-33.5,463</points>
<intersection>386 4</intersection>
<intersection>397.5 22</intersection>
<intersection>410.5 23</intersection>
<intersection>449.5 21</intersection>
<intersection>457 28</intersection>
<intersection>459 14</intersection>
<intersection>463 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-33.5,459,-19.5,459</points>
<connection>
<GID>1468</GID>
<name>K</name></connection>
<intersection>-33.5 11</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>105.5,390,109,390</points>
<connection>
<GID>1481</GID>
<name>J</name></connection>
<intersection>105.5 3</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-33.5,449.5,-32,449.5</points>
<connection>
<GID>1462</GID>
<name>IN_0</name></connection>
<intersection>-33.5 11</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-36,397.5,-33.5,397.5</points>
<connection>
<GID>1482</GID>
<name>IN_1</name></connection>
<intersection>-33.5 11</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-33.5,410.5,-25,410.5</points>
<intersection>-33.5 11</intersection>
<intersection>-25 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-25,406,-25,410.5</points>
<connection>
<GID>1470</GID>
<name>IN_1</name></connection>
<intersection>410.5 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-40,457,-33.5,457</points>
<connection>
<GID>1521</GID>
<name>OUT</name></connection>
<intersection>-33.5 11</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>105.5,415,232,415</points>
<intersection>105.5 3</intersection>
<intersection>232 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>232,384,232,415</points>
<intersection>384 33</intersection>
<intersection>415 31</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>227,384,232,384</points>
<connection>
<GID>1449</GID>
<name>J</name></connection>
<intersection>232 32</intersection></hsegment></shape></wire>
<wire>
<ID>1371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,352,108,443</points>
<intersection>352 8</intersection>
<intersection>388 1</intersection>
<intersection>443 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,388,187.5,388</points>
<connection>
<GID>1481</GID>
<name>clock</name></connection>
<connection>
<GID>1483</GID>
<name>clock</name></connection>
<connection>
<GID>1485</GID>
<name>clock</name></connection>
<connection>
<GID>1491</GID>
<name>clock</name></connection>
<connection>
<GID>1493</GID>
<name>clock</name></connection>
<intersection>108 0</intersection>
<intersection>154.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>154.5,387.5,154.5,388</points>
<connection>
<GID>1488</GID>
<name>clock</name></connection>
<intersection>388 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>108,352,200,352</points>
<connection>
<GID>1504</GID>
<name>clock</name></connection>
<connection>
<GID>1506</GID>
<name>clock</name></connection>
<connection>
<GID>1507</GID>
<name>clock</name></connection>
<connection>
<GID>1509</GID>
<name>clock</name></connection>
<connection>
<GID>1510</GID>
<name>clock</name></connection>
<connection>
<GID>1511</GID>
<name>clock</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>108,443,110.5,443</points>
<connection>
<GID>1513</GID>
<name>OUT_0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>1372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362.5,109,421.5,109</points>
<connection>
<GID>1546</GID>
<name>OUT</name></connection>
<connection>
<GID>1538</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444.5,73,444.5,109</points>
<connection>
<GID>1524</GID>
<name>IN_1</name></connection>
<intersection>109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,109,444.5,109</points>
<connection>
<GID>1538</GID>
<name>Q</name></connection>
<intersection>444.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>362,119,408.5,119</points>
<connection>
<GID>1547</GID>
<name>OUT</name></connection>
<connection>
<GID>1539</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,73,458,119</points>
<connection>
<GID>1525</GID>
<name>IN_1</name></connection>
<intersection>119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414.5,119,458,119</points>
<connection>
<GID>1539</GID>
<name>Q</name></connection>
<intersection>458 0</intersection></hsegment></shape></wire>
<wire>
<ID>1376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360.5,130,395.5,130</points>
<connection>
<GID>1548</GID>
<name>OUT</name></connection>
<connection>
<GID>1540</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>471,73,471,130</points>
<connection>
<GID>1527</GID>
<name>IN_1</name></connection>
<intersection>130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>401.5,130,471,130</points>
<connection>
<GID>1540</GID>
<name>Q</name></connection>
<intersection>471 0</intersection></hsegment></shape></wire>
<wire>
<ID>1378</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>360,139,388,139</points>
<connection>
<GID>1549</GID>
<name>OUT</name></connection>
<connection>
<GID>1541</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484,73,484,139</points>
<connection>
<GID>1528</GID>
<name>IN_1</name></connection>
<intersection>139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>394,139,484,139</points>
<connection>
<GID>1541</GID>
<name>Q</name></connection>
<intersection>484 0</intersection></hsegment></shape></wire>
<wire>
<ID>1380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,146.5,379.5,146.5</points>
<connection>
<GID>1550</GID>
<name>OUT</name></connection>
<connection>
<GID>1542</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496.5,72.5,496.5,146.5</points>
<connection>
<GID>1529</GID>
<name>IN_1</name></connection>
<intersection>146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>385.5,146.5,496.5,146.5</points>
<connection>
<GID>1542</GID>
<name>Q</name></connection>
<intersection>496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1382</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>358,154,370.5,154</points>
<connection>
<GID>1551</GID>
<name>OUT</name></connection>
<connection>
<GID>1543</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,72.5,509,154</points>
<connection>
<GID>1531</GID>
<name>IN_1</name></connection>
<intersection>154 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>376.5,154,509,154</points>
<connection>
<GID>1543</GID>
<name>Q</name></connection>
<intersection>509 0</intersection></hsegment></shape></wire>
<wire>
<ID>1384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366,107,366,158</points>
<connection>
<GID>1544</GID>
<name>OUT_0</name></connection>
<intersection>107 7</intersection>
<intersection>117 5</intersection>
<intersection>128 8</intersection>
<intersection>137 3</intersection>
<intersection>144.5 9</intersection>
<intersection>152 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>366,152,370.5,152</points>
<connection>
<GID>1543</GID>
<name>clock</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>366,137,388,137</points>
<connection>
<GID>1541</GID>
<name>clock</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>366,117,408.5,117</points>
<connection>
<GID>1539</GID>
<name>clock</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>366,107,421.5,107</points>
<connection>
<GID>1538</GID>
<name>clock</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>366,128,395.5,128</points>
<connection>
<GID>1540</GID>
<name>clock</name></connection>
<intersection>366 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>366,144.5,379.5,144.5</points>
<connection>
<GID>1542</GID>
<name>clock</name></connection>
<intersection>366 0</intersection></hsegment></shape></wire>
<wire>
<ID>1385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,103,432,158</points>
<connection>
<GID>1545</GID>
<name>OUT_0</name></connection>
<intersection>103 7</intersection>
<intersection>113 10</intersection>
<intersection>124 12</intersection>
<intersection>133 9</intersection>
<intersection>140.5 3</intersection>
<intersection>148 8</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>382.5,140.5,432,140.5</points>
<connection>
<GID>1542</GID>
<name>clear</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>424.5,103,432,103</points>
<connection>
<GID>1538</GID>
<name>clear</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>373.5,148,432,148</points>
<connection>
<GID>1543</GID>
<name>clear</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>391,133,432,133</points>
<connection>
<GID>1541</GID>
<name>clear</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>411.5,113,432,113</points>
<connection>
<GID>1539</GID>
<name>clear</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>398.5,124,432,124</points>
<connection>
<GID>1540</GID>
<name>clear</name></connection>
<intersection>432 0</intersection></hsegment></shape></wire>
<wire>
<ID>1387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534,33.5,534,36.5</points>
<intersection>33.5 2</intersection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534,36.5,539,36.5</points>
<connection>
<GID>1587</GID>
<name>IN_0</name></connection>
<intersection>534 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,33.5,534,33.5</points>
<connection>
<GID>1589</GID>
<name>OUT</name></connection>
<intersection>534 0</intersection></hsegment></shape></wire>
<wire>
<ID>1390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,388,227.5,401</points>
<intersection>388 2</intersection>
<intersection>401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220.5,401,227.5,401</points>
<connection>
<GID>1461</GID>
<name>OUT_0</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,388,227.5,388</points>
<connection>
<GID>1449</GID>
<name>K</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490,19,490,22</points>
<connection>
<GID>1489</GID>
<name>OUT</name></connection>
<intersection>19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>490,19,573,19</points>
<intersection>490 0</intersection>
<intersection>551.5 5</intersection>
<intersection>573 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>573,19,573,37.5</points>
<connection>
<GID>1595</GID>
<name>IN_0</name></connection>
<intersection>19 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>551.5,19,551.5,32</points>
<connection>
<GID>1601</GID>
<name>IN_1</name></connection>
<intersection>19 1</intersection></vsegment></shape></wire>
<wire>
<ID>1397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352.5,216.5,352.5,512.5</points>
<intersection>216.5 2</intersection>
<intersection>512.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>574,43.5,574,216.5</points>
<connection>
<GID>1595</GID>
<name>OUT</name></connection>
<intersection>216.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>352.5,216.5,574,216.5</points>
<intersection>352.5 0</intersection>
<intersection>574 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,512.5,352.5,512.5</points>
<intersection>-29 4</intersection>
<intersection>224 6</intersection>
<intersection>352.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-29,476.5,-29,512.5</points>
<intersection>476.5 5</intersection>
<intersection>512.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-33.5,476.5,-29,476.5</points>
<connection>
<GID>1496</GID>
<name>IN_0</name></connection>
<intersection>-29 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>224,390,224,512.5</points>
<connection>
<GID>1449</GID>
<name>clear</name></connection>
<intersection>512.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>548,34,548,35.5</points>
<intersection>34 2</intersection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>545,35.5,548,35.5</points>
<connection>
<GID>1587</GID>
<name>OUT</name></connection>
<intersection>548 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>548,34,551.5,34</points>
<connection>
<GID>1601</GID>
<name>IN_0</name></connection>
<intersection>548 0</intersection></hsegment></shape></wire>
<wire>
<ID>1399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>575,33,575,37.5</points>
<connection>
<GID>1595</GID>
<name>IN_1</name></connection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>557.5,33,575,33</points>
<connection>
<GID>1601</GID>
<name>OUT</name></connection>
<intersection>575 0</intersection></hsegment></shape></wire>
<wire>
<ID>1407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,384,216,385</points>
<intersection>384 2</intersection>
<intersection>385 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,385,216,385</points>
<connection>
<GID>1460</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,384,221,384</points>
<connection>
<GID>1449</GID>
<name>Q</name></connection>
<intersection>216 0</intersection></hsegment></shape></wire>
<wire>
<ID>1408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,388,166.5,471</points>
<intersection>388 2</intersection>
<intersection>471 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,471,166.5,471</points>
<connection>
<GID>1456</GID>
<name>IN_0</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,388,221,388</points>
<connection>
<GID>1449</GID>
<name>nQ</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,458,-44,479.5</points>
<connection>
<GID>1479</GID>
<name>OUT_0</name></connection>
<intersection>458 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,458,-44,458</points>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>1229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,16,326,167.5</points>
<connection>
<GID>1472</GID>
<name>OUT_0</name></connection>
<intersection>16 13</intersection>
<intersection>110 1</intersection>
<intersection>120 3</intersection>
<intersection>131 5</intersection>
<intersection>140 7</intersection>
<intersection>147.5 9</intersection>
<intersection>155 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326,110,356.5,110</points>
<connection>
<GID>1546</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>326,120,356,120</points>
<connection>
<GID>1547</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>326,131,354.5,131</points>
<connection>
<GID>1548</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>326,140,354,140</points>
<connection>
<GID>1549</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>326,147.5,353,147.5</points>
<connection>
<GID>1550</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>326,155,352,155</points>
<connection>
<GID>1551</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>326,16,539,16</points>
<intersection>326 0</intersection>
<intersection>539 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>539,16,539,34.5</points>
<connection>
<GID>1587</GID>
<name>IN_1</name></connection>
<intersection>16 13</intersection></vsegment></shape></wire>
<wire>
<ID>1230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,63.5,445.5,67</points>
<connection>
<GID>1524</GID>
<name>OUT</name></connection>
<intersection>63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,63.5,446.5,63.5</points>
<connection>
<GID>1566</GID>
<name>IN_0</name></connection>
<intersection>445.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,63,459,67</points>
<connection>
<GID>1525</GID>
<name>OUT</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459,63,462.5,63</points>
<connection>
<GID>1414</GID>
<name>IN_0</name></connection>
<intersection>459 0</intersection></hsegment></shape></wire>
<wire>
<ID>1232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>472,63,472,67</points>
<connection>
<GID>1527</GID>
<name>OUT</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>472,63,476,63</points>
<connection>
<GID>1423</GID>
<name>IN_0</name></connection>
<intersection>472 0</intersection></hsegment></shape></wire>
<wire>
<ID>1233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488,63,488,67</points>
<intersection>63 1</intersection>
<intersection>67 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>488,63,491,63</points>
<connection>
<GID>1430</GID>
<name>IN_0</name></connection>
<intersection>488 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>485,67,488,67</points>
<connection>
<GID>1528</GID>
<name>OUT</name></connection>
<intersection>488 0</intersection></hsegment></shape></wire>
<wire>
<ID>1234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497.5,64.5,497.5,66.5</points>
<connection>
<GID>1529</GID>
<name>OUT</name></connection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,64.5,501.5,64.5</points>
<intersection>497.5 0</intersection>
<intersection>501.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>501.5,63,501.5,64.5</points>
<connection>
<GID>1435</GID>
<name>IN_0</name></connection>
<intersection>64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,64.5,510,66.5</points>
<connection>
<GID>1531</GID>
<name>OUT</name></connection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,64.5,514.5,64.5</points>
<intersection>510 0</intersection>
<intersection>514.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>514.5,63,514.5,64.5</points>
<connection>
<GID>1441</GID>
<name>IN_0</name></connection>
<intersection>64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,55.5,456.5,63.5</points>
<connection>
<GID>1445</GID>
<name>IN_0</name></connection>
<intersection>63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,63.5,456.5,63.5</points>
<connection>
<GID>1566</GID>
<name>OUT_0</name></connection>
<intersection>456.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>471.5,55.5,471.5,63</points>
<connection>
<GID>1448</GID>
<name>IN_0</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>468.5,63,471.5,63</points>
<connection>
<GID>1414</GID>
<name>OUT_0</name></connection>
<intersection>471.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>486.5,55.5,486.5,63</points>
<connection>
<GID>1451</GID>
<name>IN_0</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>482,63,486.5,63</points>
<connection>
<GID>1423</GID>
<name>OUT_0</name></connection>
<intersection>486.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498,56,498,63</points>
<connection>
<GID>1453</GID>
<name>IN_0</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497,63,498,63</points>
<connection>
<GID>1430</GID>
<name>OUT_0</name></connection>
<intersection>498 0</intersection></hsegment></shape></wire>
<wire>
<ID>1240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,55.5,511,63</points>
<connection>
<GID>1455</GID>
<name>IN_0</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507.5,63,511,63</points>
<connection>
<GID>1435</GID>
<name>OUT_0</name></connection>
<intersection>511 0</intersection></hsegment></shape></wire>
<wire>
<ID>1241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524,56,524,63</points>
<connection>
<GID>1458</GID>
<name>IN_0</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>520.5,63,524,63</points>
<connection>
<GID>1441</GID>
<name>OUT_0</name></connection>
<intersection>524 0</intersection></hsegment></shape></wire>
<wire>
<ID>1242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,46,456.5,51.5</points>
<connection>
<GID>1445</GID>
<name>OUT_0</name></connection>
<intersection>46 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>471.5,40,471.5,46</points>
<connection>
<GID>1475</GID>
<name>IN_3</name></connection>
<intersection>46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>456.5,46,471.5,46</points>
<intersection>456.5 0</intersection>
<intersection>471.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>471.5,46.5,471.5,51.5</points>
<connection>
<GID>1448</GID>
<name>OUT_0</name></connection>
<intersection>46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>473.5,40,473.5,46.5</points>
<connection>
<GID>1475</GID>
<name>IN_2</name></connection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>471.5,46.5,473.5,46.5</points>
<intersection>471.5 0</intersection>
<intersection>473.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>486.5,46,486.5,51.5</points>
<connection>
<GID>1451</GID>
<name>OUT_0</name></connection>
<intersection>46 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>475.5,40,475.5,46</points>
<connection>
<GID>1475</GID>
<name>IN_1</name></connection>
<intersection>46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>475.5,46,486.5,46</points>
<intersection>475.5 1</intersection>
<intersection>486.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498,45,498,52</points>
<connection>
<GID>1453</GID>
<name>OUT_0</name></connection>
<intersection>45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>477.5,40,477.5,45</points>
<connection>
<GID>1475</GID>
<name>IN_0</name></connection>
<intersection>45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>477.5,45,498,45</points>
<intersection>477.5 1</intersection>
<intersection>498 0</intersection></hsegment></shape></wire>
<wire>
<ID>1246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,46.5,511,51.5</points>
<connection>
<GID>1455</GID>
<name>OUT_0</name></connection>
<intersection>46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>510,41,510,46.5</points>
<connection>
<GID>1486</GID>
<name>IN_1</name></connection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>510,46.5,511,46.5</points>
<intersection>510 1</intersection>
<intersection>511 0</intersection></hsegment></shape></wire>
<wire>
<ID>1247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524,46.5,524,52</points>
<connection>
<GID>1458</GID>
<name>OUT_0</name></connection>
<intersection>46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>512,41,512,46.5</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>512,46.5,524,46.5</points>
<intersection>512 1</intersection>
<intersection>524 0</intersection></hsegment></shape></wire>
<wire>
<ID>1248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>474.5,31,474.5,34</points>
<connection>
<GID>1475</GID>
<name>OUT</name></connection>
<intersection>31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>489,28,489,31</points>
<connection>
<GID>1489</GID>
<name>IN_1</name></connection>
<intersection>29.5 3</intersection>
<intersection>31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>474.5,31,489,31</points>
<intersection>474.5 0</intersection>
<intersection>489 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>489,29.5,523,29.5</points>
<intersection>489 1</intersection>
<intersection>523 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>523,29.5,523,32.5</points>
<connection>
<GID>1589</GID>
<name>IN_1</name></connection>
<intersection>29.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,31.5,511,35</points>
<connection>
<GID>1486</GID>
<name>OUT</name></connection>
<intersection>31.5 2</intersection>
<intersection>34.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>491,28,491,31.5</points>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>491,31.5,511,31.5</points>
<intersection>491 1</intersection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>511,34.5,523,34.5</points>
<connection>
<GID>1589</GID>
<name>IN_0</name></connection>
<intersection>511 0</intersection></hsegment></shape></wire>
<wire>
<ID>1253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-109.5,292,-102,292</points>
<connection>
<GID>1523</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1522</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,290,-52,290</points>
<connection>
<GID>1533</GID>
<name>IN_0</name></connection>
<connection>
<GID>1553</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,281.5,-56,287</points>
<intersection>281.5 2</intersection>
<intersection>287 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,287,-52,287</points>
<connection>
<GID>1533</GID>
<name>clock</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-102,281.5,-56,281.5</points>
<intersection>-102 3</intersection>
<intersection>-60 4</intersection>
<intersection>-56 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-102,281.5,-102,289</points>
<connection>
<GID>1522</GID>
<name>clock</name></connection>
<intersection>281.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-60,281.5,-60,284.5</points>
<connection>
<GID>1534</GID>
<name>CLK</name></connection>
<intersection>281.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81.5,278,-81.5,298</points>
<connection>
<GID>1526</GID>
<name>IN_1</name></connection>
<intersection>278 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81.5,278,-46,278</points>
<intersection>-81.5 0</intersection>
<intersection>-46 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-46,278,-46,287</points>
<connection>
<GID>1533</GID>
<name>OUTINV_0</name></connection>
<intersection>278 1</intersection></vsegment></shape></wire>
<wire>
<ID>1257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83.5,292,-83.5,298</points>
<connection>
<GID>1526</GID>
<name>IN_0</name></connection>
<intersection>292 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-96,292,-83.5,292</points>
<connection>
<GID>1522</GID>
<name>OUT_0</name></connection>
<intersection>-83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82.5,304,-82.5,456</points>
<connection>
<GID>1526</GID>
<name>OUT</name></connection>
<intersection>456 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82.5,456,-46,456</points>
<connection>
<GID>1521</GID>
<name>IN_1</name></connection>
<intersection>-82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-96,289,-90.5,289</points>
<connection>
<GID>1522</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>1530</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,249,-49,284</points>
<connection>
<GID>1533</GID>
<name>clear</name></connection>
<intersection>249 3</intersection>
<intersection>276.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-86.5,276.5,-49,276.5</points>
<intersection>-86.5 2</intersection>
<intersection>-49 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-86.5,276.5,-86.5,289</points>
<connection>
<GID>1530</GID>
<name>OUT_0</name></connection>
<intersection>276.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-49,249,-33.5,249</points>
<connection>
<GID>1585</GID>
<name>clear</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>1261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,231.5,255,287</points>
<intersection>231.5 2</intersection>
<intersection>287 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,287,255,287</points>
<connection>
<GID>1555</GID>
<name>OUT</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,231.5,255,231.5</points>
<intersection>30 15</intersection>
<intersection>79.5 14</intersection>
<intersection>105.5 10</intersection>
<intersection>135.5 18</intersection>
<intersection>174 16</intersection>
<intersection>222.5 17</intersection>
<intersection>255 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>105.5,231.5,105.5,257.5</points>
<connection>
<GID>1560</GID>
<name>clear</name></connection>
<intersection>231.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>79.5,231.5,79.5,257</points>
<connection>
<GID>1558</GID>
<name>clear</name></connection>
<intersection>231.5 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>30,231.5,30,257.5</points>
<connection>
<GID>1557</GID>
<name>clear</name></connection>
<intersection>231.5 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>174,231.5,174,255</points>
<connection>
<GID>1562</GID>
<name>clear</name></connection>
<intersection>231.5 2</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>222.5,231.5,222.5,254.5</points>
<connection>
<GID>1563</GID>
<name>clear</name></connection>
<intersection>231.5 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>135.5,231.5,135.5,257</points>
<connection>
<GID>1561</GID>
<name>clear</name></connection>
<intersection>231.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,219,39,269.5</points>
<intersection>219 8</intersection>
<intersection>225 5</intersection>
<intersection>234.5 3</intersection>
<intersection>263.5 2</intersection>
<intersection>269.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,269.5,43.5,269.5</points>
<connection>
<GID>1565</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,263.5,39,263.5</points>
<connection>
<GID>1557</GID>
<name>Q</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,234.5,242,234.5</points>
<connection>
<GID>1584</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>39,225,58,225</points>
<intersection>39 0</intersection>
<intersection>58 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>58,192.5,58,225</points>
<connection>
<GID>1431</GID>
<name>IN_0</name></connection>
<intersection>225 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>39,219,45,219</points>
<connection>
<GID>1556</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>1263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,254,35,259.5</points>
<intersection>254 3</intersection>
<intersection>259.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,259.5,35,259.5</points>
<connection>
<GID>1557</GID>
<name>nQ</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,254,42.5,254</points>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>1264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,262,53.5,271.5</points>
<intersection>262 1</intersection>
<intersection>270.5 2</intersection>
<intersection>271.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,262,57.5,262</points>
<connection>
<GID>1577</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,270.5,53.5,270.5</points>
<connection>
<GID>1565</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53.5,271.5,84.5,271.5</points>
<connection>
<GID>1568</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,251,54,260</points>
<intersection>251 2</intersection>
<intersection>253 3</intersection>
<intersection>260 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,260,57.5,260</points>
<connection>
<GID>1577</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,251,87,251</points>
<connection>
<GID>1569</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>48.5,253,54,253</points>
<connection>
<GID>1567</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>1266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,193,83.5,269.5</points>
<intersection>193 9</intersection>
<intersection>219.5 5</intersection>
<intersection>235.5 3</intersection>
<intersection>263 2</intersection>
<intersection>269.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,269.5,84.5,269.5</points>
<connection>
<GID>1568</GID>
<name>IN_1</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,263,83.5,263</points>
<connection>
<GID>1558</GID>
<name>Q</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83.5,235.5,242,235.5</points>
<connection>
<GID>1584</GID>
<name>IN_1</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>83.5,219.5,88,219.5</points>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>70.5,193,83.5,193</points>
<intersection>70.5 10</intersection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>70.5,191.5,70.5,193</points>
<connection>
<GID>1432</GID>
<name>IN_0</name></connection>
<intersection>193 9</intersection></vsegment></shape></wire>
<wire>
<ID>1267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,107.5,54,219</points>
<intersection>107.5 5</intersection>
<intersection>204 10</intersection>
<intersection>219 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,219,54,219</points>
<connection>
<GID>1556</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54,107.5,356.5,107.5</points>
<intersection>54 0</intersection>
<intersection>356.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>356.5,107.5,356.5,108</points>
<connection>
<GID>1546</GID>
<name>IN_1</name></connection>
<intersection>107.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>54,204,261.5,204</points>
<connection>
<GID>1410</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>1268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,270,92,270.5</points>
<intersection>270 2</intersection>
<intersection>270.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,270.5,92,270.5</points>
<connection>
<GID>1568</GID>
<name>OUT</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,270,114,270</points>
<connection>
<GID>1570</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection>
<intersection>94 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>94,263,94,270</points>
<connection>
<GID>1579</GID>
<name>IN_0</name></connection>
<intersection>270 2</intersection></vsegment></shape></wire>
<wire>
<ID>1269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,253,85,259</points>
<intersection>253 2</intersection>
<intersection>259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,259,85,259</points>
<connection>
<GID>1558</GID>
<name>nQ</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,253,87,253</points>
<connection>
<GID>1569</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>1270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,249.5,93.5,261</points>
<intersection>249.5 3</intersection>
<intersection>252 1</intersection>
<intersection>261 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,252,93.5,252</points>
<connection>
<GID>1569</GID>
<name>OUT</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,261,94,261</points>
<connection>
<GID>1579</GID>
<name>IN_1</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>93.5,249.5,116.5,249.5</points>
<connection>
<GID>1571</GID>
<name>IN_1</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,192.5,110.5,290</points>
<intersection>192.5 13</intersection>
<intersection>219.5 9</intersection>
<intersection>236.5 2</intersection>
<intersection>263.5 1</intersection>
<intersection>268 5</intersection>
<intersection>290 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,263.5,110.5,263.5</points>
<connection>
<GID>1560</GID>
<name>Q</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,236.5,242,236.5</points>
<connection>
<GID>1584</GID>
<name>IN_2</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>110.5,268,114,268</points>
<connection>
<GID>1570</GID>
<name>IN_1</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>110.5,290,244,290</points>
<connection>
<GID>1555</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>110.5,219.5,117.5,219.5</points>
<connection>
<GID>1564</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>110.5,192.5,134.5,192.5</points>
<connection>
<GID>1433</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1272</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,269,140.5,269</points>
<connection>
<GID>1570</GID>
<name>OUT</name></connection>
<connection>
<GID>1572</GID>
<name>IN_0</name></connection>
<intersection>122.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122.5,262.5,122.5,269</points>
<connection>
<GID>1580</GID>
<name>IN_0</name></connection>
<intersection>269 1</intersection></vsegment></shape></wire>
<wire>
<ID>1273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,249.5,122.5,260.5</points>
<connection>
<GID>1580</GID>
<name>IN_1</name></connection>
<connection>
<GID>1571</GID>
<name>OUT</name></connection>
<intersection>249.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,249.5,142,249.5</points>
<connection>
<GID>1573</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,251.5,112,259.5</points>
<intersection>251.5 2</intersection>
<intersection>259.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,259.5,112,259.5</points>
<connection>
<GID>1560</GID>
<name>nQ</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112,251.5,116.5,251.5</points>
<connection>
<GID>1571</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>1275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,219.5,138.5,288</points>
<connection>
<GID>1561</GID>
<name>Q</name></connection>
<intersection>219.5 10</intersection>
<intersection>237.5 2</intersection>
<intersection>267 6</intersection>
<intersection>288 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138.5,237.5,242,237.5</points>
<connection>
<GID>1584</GID>
<name>IN_3</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>138.5,267,140.5,267</points>
<connection>
<GID>1572</GID>
<name>IN_1</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>138.5,288,244,288</points>
<connection>
<GID>1555</GID>
<name>IN_1</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>138.5,219.5,146,219.5</points>
<connection>
<GID>1576</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection>
<intersection>141.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>141.5,192.5,141.5,219.5</points>
<connection>
<GID>1434</GID>
<name>IN_0</name></connection>
<intersection>219.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>1276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,251.5,139.5,259</points>
<intersection>251.5 2</intersection>
<intersection>259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,259,139.5,259</points>
<connection>
<GID>1561</GID>
<name>nQ</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,251.5,142,251.5</points>
<connection>
<GID>1573</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,262,149.5,270</points>
<intersection>262 2</intersection>
<intersection>268 1</intersection>
<intersection>270 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146.5,268,149.5,268</points>
<connection>
<GID>1572</GID>
<name>OUT</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149.5,262,151.5,262</points>
<connection>
<GID>1581</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>149.5,270,187.5,270</points>
<connection>
<GID>1574</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,250.5,150,260</points>
<intersection>250.5 1</intersection>
<intersection>260 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,250.5,188,250.5</points>
<connection>
<GID>1573</GID>
<name>OUT</name></connection>
<connection>
<GID>1575</GID>
<name>IN_1</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>150,260,151.5,260</points>
<connection>
<GID>1581</GID>
<name>IN_1</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>1279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,193,182,286</points>
<intersection>193 14</intersection>
<intersection>219.5 9</intersection>
<intersection>238.5 3</intersection>
<intersection>261 1</intersection>
<intersection>268 10</intersection>
<intersection>286 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,261,182,261</points>
<connection>
<GID>1562</GID>
<name>Q</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>182,238.5,242,238.5</points>
<connection>
<GID>1584</GID>
<name>IN_4</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182,286,244,286</points>
<connection>
<GID>1555</GID>
<name>IN_2</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>182,219.5,192,219.5</points>
<connection>
<GID>1578</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>182,268,187.5,268</points>
<connection>
<GID>1574</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>182,193,199,193</points>
<connection>
<GID>1436</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>1280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,252.5,179.5,257</points>
<intersection>252.5 2</intersection>
<intersection>257 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,257,179.5,257</points>
<connection>
<GID>1562</GID>
<name>nQ</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179.5,252.5,188,252.5</points>
<connection>
<GID>1575</GID>
<name>IN_0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,261.5,194.5,269</points>
<intersection>261.5 2</intersection>
<intersection>269 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,269,194.5,269</points>
<connection>
<GID>1574</GID>
<name>OUT</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,261.5,195.5,261.5</points>
<connection>
<GID>1582</GID>
<name>IN_0</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,251.5,194.5,259.5</points>
<intersection>251.5 1</intersection>
<intersection>259.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,251.5,194.5,251.5</points>
<connection>
<GID>1575</GID>
<name>OUT</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,259.5,195.5,259.5</points>
<connection>
<GID>1582</GID>
<name>IN_1</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,242,219.5,242</points>
<intersection>1.5 16</intersection>
<intersection>19 13</intersection>
<intersection>76 12</intersection>
<intersection>101.5 6</intersection>
<intersection>129.5 7</intersection>
<intersection>167.5 11</intersection>
<intersection>219.5 28</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>101.5,242,101.5,261.5</points>
<intersection>242 1</intersection>
<intersection>261.5 19</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>129.5,242,129.5,261</points>
<intersection>242 1</intersection>
<intersection>261 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>167.5,242,167.5,259</points>
<intersection>242 1</intersection>
<intersection>259 18</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>76,242,76,261</points>
<intersection>242 1</intersection>
<intersection>261 22</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>19,242,19,261.5</points>
<intersection>242 1</intersection>
<intersection>261.5 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>129.5,261,132.5,261</points>
<connection>
<GID>1561</GID>
<name>clock</name></connection>
<intersection>129.5 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>19,261.5,27,261.5</points>
<connection>
<GID>1557</GID>
<name>clock</name></connection>
<intersection>19 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>1.5,212.5,1.5,242</points>
<intersection>212.5 17</intersection>
<intersection>241.5 37</intersection>
<intersection>242 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>1.5,212.5,240,212.5</points>
<intersection>1.5 16</intersection>
<intersection>45 34</intersection>
<intersection>88 25</intersection>
<intersection>117.5 26</intersection>
<intersection>146 24</intersection>
<intersection>191 23</intersection>
<intersection>240 35</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>167.5,259,171,259</points>
<connection>
<GID>1562</GID>
<name>clock</name></connection>
<intersection>167.5 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>101.5,261.5,102.5,261.5</points>
<connection>
<GID>1560</GID>
<name>clock</name></connection>
<intersection>101.5 6</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>76,261,76.5,261</points>
<connection>
<GID>1558</GID>
<name>clock</name></connection>
<intersection>76 12</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>191,212.5,191,216.5</points>
<intersection>212.5 17</intersection>
<intersection>216.5 36</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>146,212.5,146,216.5</points>
<connection>
<GID>1576</GID>
<name>clock</name></connection>
<intersection>212.5 17</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>88,212.5,88,216.5</points>
<connection>
<GID>1559</GID>
<name>clock</name></connection>
<intersection>212.5 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>117.5,212.5,117.5,216.5</points>
<connection>
<GID>1564</GID>
<name>clock</name></connection>
<intersection>212.5 17</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>219.5,242,219.5,258.5</points>
<connection>
<GID>1563</GID>
<name>clock</name></connection>
<intersection>242 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>45,212.5,45,216</points>
<connection>
<GID>1556</GID>
<name>clock</name></connection>
<intersection>212.5 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>240,212.5,240,216</points>
<connection>
<GID>1583</GID>
<name>clock</name></connection>
<intersection>212.5 17</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>191,216.5,192,216.5</points>
<connection>
<GID>1578</GID>
<name>clock</name></connection>
<intersection>191 23</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-39.5,241.5,1.5,241.5</points>
<connection>
<GID>1413</GID>
<name>OUT</name></connection>
<intersection>-37 38</intersection>
<intersection>1.5 16</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>-37,241.5,-37,252</points>
<intersection>241.5 37</intersection>
<intersection>252 39</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-37,252,-36.5,252</points>
<connection>
<GID>1585</GID>
<name>clock</name></connection>
<intersection>-37 38</intersection></hsegment></shape></wire>
<wire>
<ID>1284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,193.5,234.5,284</points>
<intersection>193.5 9</intersection>
<intersection>219 13</intersection>
<intersection>239.5 2</intersection>
<intersection>260.5 11</intersection>
<intersection>284 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>234.5,239.5,242,239.5</points>
<connection>
<GID>1584</GID>
<name>IN_5</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>234.5,284,244,284</points>
<connection>
<GID>1555</GID>
<name>IN_3</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>204.5,193.5,234.5,193.5</points>
<connection>
<GID>1437</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>225.5,260.5,234.5,260.5</points>
<connection>
<GID>1563</GID>
<name>Q</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>234.5,219,240,219</points>
<connection>
<GID>1583</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1285</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>95.5,118,95.5,219.5</points>
<intersection>118 11</intersection>
<intersection>205 14</intersection>
<intersection>219.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94,219.5,95.5,219.5</points>
<connection>
<GID>1559</GID>
<name>OUT_0</name></connection>
<intersection>95.5 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>95.5,118,356,118</points>
<connection>
<GID>1547</GID>
<name>IN_1</name></connection>
<intersection>95.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>95.5,205,261.5,205</points>
<connection>
<GID>1410</GID>
<name>IN_1</name></connection>
<intersection>95.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1286</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>125,129,125,219.5</points>
<intersection>129 7</intersection>
<intersection>206 12</intersection>
<intersection>219.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>123.5,219.5,125,219.5</points>
<connection>
<GID>1564</GID>
<name>OUT_0</name></connection>
<intersection>125 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125,129,354.5,129</points>
<connection>
<GID>1548</GID>
<name>IN_1</name></connection>
<intersection>125 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>125,206,261.5,206</points>
<connection>
<GID>1410</GID>
<name>IN_2</name></connection>
<intersection>125 3</intersection></hsegment></shape></wire>
<wire>
<ID>1287</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>152,138,152,219.5</points>
<connection>
<GID>1576</GID>
<name>OUT_0</name></connection>
<intersection>138 7</intersection>
<intersection>207 15</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>152,138,354,138</points>
<connection>
<GID>1549</GID>
<name>IN_1</name></connection>
<intersection>152 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>152,207,261.5,207</points>
<connection>
<GID>1410</GID>
<name>IN_3</name></connection>
<intersection>152 3</intersection></hsegment></shape></wire>
<wire>
<ID>1288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,145.5,210,219.5</points>
<intersection>145.5 5</intersection>
<intersection>208 10</intersection>
<intersection>219.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,219.5,210,219.5</points>
<connection>
<GID>1578</GID>
<name>OUT_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>210,145.5,353,145.5</points>
<connection>
<GID>1550</GID>
<name>IN_1</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>210,208,261.5,208</points>
<connection>
<GID>1410</GID>
<name>IN_4</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>1289</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>253,153,253,219</points>
<intersection>153 10</intersection>
<intersection>209 16</intersection>
<intersection>219 13</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>253,153,352,153</points>
<connection>
<GID>1551</GID>
<name>IN_1</name></connection>
<intersection>253 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>246,219,253,219</points>
<connection>
<GID>1583</GID>
<name>OUT_0</name></connection>
<intersection>253 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>253,209,261.5,209</points>
<connection>
<GID>1410</GID>
<name>IN_5</name></connection>
<intersection>253 3</intersection></hsegment></shape></wire>
<wire>
<ID>1290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,263.5,24,276</points>
<intersection>263.5 8</intersection>
<intersection>276 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>15.5,276,24,276</points>
<intersection>15.5 9</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>24,263.5,27,263.5</points>
<connection>
<GID>1557</GID>
<name>J</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>15.5,275.5,15.5,287.5</points>
<connection>
<GID>1422</GID>
<name>IN_0</name></connection>
<intersection>276 6</intersection>
<intersection>287.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-25.5,287.5,15.5,287.5</points>
<intersection>-25.5 14</intersection>
<intersection>15.5 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-25.5,284,-25.5,287.5</points>
<intersection>284 15</intersection>
<intersection>287.5 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-36,284,-25.5,284</points>
<connection>
<GID>1439</GID>
<name>OUT</name></connection>
<intersection>-25.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>1291</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>9,283,207,283</points>
<intersection>9 7</intersection>
<intersection>64.5 6</intersection>
<intersection>101 10</intersection>
<intersection>129.5 12</intersection>
<intersection>159.5 14</intersection>
<intersection>207 16</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>64.5,278,64.5,283</points>
<connection>
<GID>1424</GID>
<name>IN_1</name></connection>
<intersection>283 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>9,276,9,283</points>
<intersection>276 20</intersection>
<intersection>283 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>101,278.5,101,283</points>
<connection>
<GID>1425</GID>
<name>IN_1</name></connection>
<intersection>283 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>129.5,278,129.5,283</points>
<connection>
<GID>1426</GID>
<name>IN_1</name></connection>
<intersection>283 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>159.5,278,159.5,283</points>
<connection>
<GID>1427</GID>
<name>IN_1</name></connection>
<intersection>283 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>207,280,207,283</points>
<connection>
<GID>1428</GID>
<name>IN_1</name></connection>
<intersection>283 4</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-21.5,276,13.5,276</points>
<intersection>-21.5 23</intersection>
<intersection>9 7</intersection>
<intersection>13.5 26</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-21.5,140.5,-21.5,276</points>
<intersection>140.5 24</intersection>
<intersection>276 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-21.5,140.5,42.5,140.5</points>
<intersection>-21.5 23</intersection>
<intersection>42.5 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>42.5,140.5,42.5,141.5</points>
<connection>
<GID>1429</GID>
<name>OUT</name></connection>
<intersection>140.5 24</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>13.5,275.5,13.5,276</points>
<connection>
<GID>1422</GID>
<name>IN_1</name></connection>
<intersection>276 20</intersection></vsegment></shape></wire>
<wire>
<ID>1292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,259.5,14.5,269.5</points>
<connection>
<GID>1422</GID>
<name>OUT</name></connection>
<intersection>259.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,259.5,27,259.5</points>
<connection>
<GID>1557</GID>
<name>K</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,169.5,63,181</points>
<connection>
<GID>1416</GID>
<name>IN_1</name></connection>
<intersection>181 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58,181,58,186.5</points>
<connection>
<GID>1431</GID>
<name>OUT_0</name></connection>
<intersection>181 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58,181,63,181</points>
<intersection>58 1</intersection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>1294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,169.5,65,181</points>
<connection>
<GID>1416</GID>
<name>IN_0</name></connection>
<intersection>181 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70.5,181,70.5,185.5</points>
<connection>
<GID>1432</GID>
<name>OUT_0</name></connection>
<intersection>181 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>65,181,70.5,181</points>
<intersection>65 0</intersection>
<intersection>70.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,147.5,41.5,160</points>
<connection>
<GID>1429</GID>
<name>IN_2</name></connection>
<intersection>160 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64,160,64,163.5</points>
<connection>
<GID>1416</GID>
<name>OUT</name></connection>
<intersection>160 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41.5,160,64,160</points>
<intersection>41.5 0</intersection>
<intersection>64 1</intersection></hsegment></shape></wire>
<wire>
<ID>1296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,183,139,185</points>
<connection>
<GID>1419</GID>
<name>IN_0</name></connection>
<intersection>185 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>141.5,185,141.5,186.5</points>
<connection>
<GID>1434</GID>
<name>OUT_0</name></connection>
<intersection>185 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>139,185,141.5,185</points>
<intersection>139 0</intersection>
<intersection>141.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,183,137,185</points>
<connection>
<GID>1419</GID>
<name>IN_1</name></connection>
<intersection>185 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>134.5,185,134.5,186.5</points>
<connection>
<GID>1433</GID>
<name>OUT_0</name></connection>
<intersection>185 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134.5,185,137,185</points>
<intersection>134.5 1</intersection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>1298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,147.5,43.5,158</points>
<connection>
<GID>1429</GID>
<name>IN_1</name></connection>
<intersection>158 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>138,158,138,177</points>
<connection>
<GID>1419</GID>
<name>OUT</name></connection>
<intersection>158 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>43.5,158,138,158</points>
<intersection>43.5 0</intersection>
<intersection>138 1</intersection></hsegment></shape></wire>
<wire>
<ID>1299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202,184.5,202,186</points>
<connection>
<GID>1421</GID>
<name>IN_0</name></connection>
<intersection>186 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>204.5,186,204.5,187.5</points>
<connection>
<GID>1437</GID>
<name>OUT_0</name></connection>
<intersection>186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>202,186,204.5,186</points>
<intersection>202 0</intersection>
<intersection>204.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200,184.5,200,186</points>
<connection>
<GID>1421</GID>
<name>IN_1</name></connection>
<intersection>186 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>199,186,199,187</points>
<connection>
<GID>1436</GID>
<name>OUT_0</name></connection>
<intersection>186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>199,186,200,186</points>
<intersection>199 1</intersection>
<intersection>200 0</intersection></hsegment></shape></wire>
<wire>
<ID>1301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,147.5,45.5,155.5</points>
<connection>
<GID>1429</GID>
<name>IN_0</name></connection>
<intersection>155.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>201,155.5,201,178.5</points>
<connection>
<GID>1421</GID>
<name>OUT</name></connection>
<intersection>155.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,155.5,201,155.5</points>
<intersection>45.5 0</intersection>
<intersection>201 1</intersection></hsegment></shape></wire>
<wire>
<ID>1302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,261,74,278.5</points>
<intersection>261 2</intersection>
<intersection>263 1</intersection>
<intersection>278.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,263,76.5,263</points>
<connection>
<GID>1558</GID>
<name>J</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,261,74,261</points>
<connection>
<GID>1577</GID>
<name>OUT</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>66.5,278.5,74,278.5</points>
<intersection>66.5 4</intersection>
<intersection>74 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>66.5,278,66.5,278.5</points>
<connection>
<GID>1424</GID>
<name>IN_0</name></connection>
<intersection>278.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,259,65.5,272</points>
<connection>
<GID>1424</GID>
<name>OUT</name></connection>
<intersection>259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,259,76.5,259</points>
<connection>
<GID>1558</GID>
<name>K</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,263.5,102,272.5</points>
<connection>
<GID>1425</GID>
<name>OUT</name></connection>
<intersection>263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,263.5,102.5,263.5</points>
<connection>
<GID>1560</GID>
<name>J</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>1305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,271,109.5,278.5</points>
<intersection>271 1</intersection>
<intersection>278.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,271,109.5,271</points>
<intersection>100 4</intersection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,278.5,109.5,278.5</points>
<connection>
<GID>1425</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,259.5,100,271</points>
<connection>
<GID>1579</GID>
<name>OUT</name></connection>
<intersection>259.5 6</intersection>
<intersection>271 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>100,259.5,102.5,259.5</points>
<connection>
<GID>1560</GID>
<name>K</name></connection>
<intersection>100 4</intersection></hsegment></shape></wire>
<wire>
<ID>1306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128.5,270.5,135,270.5</points>
<intersection>128.5 3</intersection>
<intersection>135 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,261.5,128.5,270.5</points>
<connection>
<GID>1580</GID>
<name>OUT</name></connection>
<intersection>263 7</intersection>
<intersection>270.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>135,270.5,135,278</points>
<intersection>270.5 1</intersection>
<intersection>278 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>131.5,278,135,278</points>
<connection>
<GID>1426</GID>
<name>IN_0</name></connection>
<intersection>135 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>128.5,263,132.5,263</points>
<connection>
<GID>1561</GID>
<name>J</name></connection>
<intersection>128.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,259,130.5,272</points>
<connection>
<GID>1426</GID>
<name>OUT</name></connection>
<intersection>259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,259,132.5,259</points>
<connection>
<GID>1561</GID>
<name>K</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157.5,261,171,261</points>
<connection>
<GID>1581</GID>
<name>OUT</name></connection>
<connection>
<GID>1562</GID>
<name>J</name></connection>
<intersection>164.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>164.5,261,164.5,279</points>
<intersection>261 1</intersection>
<intersection>279 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>161.5,279,164.5,279</points>
<intersection>161.5 6</intersection>
<intersection>164.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>161.5,278,161.5,279</points>
<connection>
<GID>1427</GID>
<name>IN_0</name></connection>
<intersection>279 5</intersection></vsegment></shape></wire>
<wire>
<ID>1309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,257,160.5,272</points>
<connection>
<GID>1427</GID>
<name>OUT</name></connection>
<intersection>257 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,257,171,257</points>
<connection>
<GID>1562</GID>
<name>K</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201.5,260.5,219.5,260.5</points>
<connection>
<GID>1582</GID>
<name>OUT</name></connection>
<connection>
<GID>1563</GID>
<name>J</name></connection>
<intersection>210 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>210,260.5,210,281.5</points>
<intersection>260.5 1</intersection>
<intersection>281.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>209,281.5,210,281.5</points>
<intersection>209 15</intersection>
<intersection>210 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>209,280,209,281.5</points>
<connection>
<GID>1428</GID>
<name>IN_0</name></connection>
<intersection>281.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>1311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,256.5,208,274</points>
<connection>
<GID>1428</GID>
<name>OUT</name></connection>
<intersection>256.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,256.5,219.5,256.5</points>
<connection>
<GID>1563</GID>
<name>K</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>1312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,290,-37,290</points>
<connection>
<GID>1439</GID>
<name>IN_1</name></connection>
<connection>
<GID>1533</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,290,-35,291</points>
<connection>
<GID>1439</GID>
<name>IN_0</name></connection>
<intersection>291 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-29,291,-29,292.5</points>
<connection>
<GID>1412</GID>
<name>OUT_0</name></connection>
<intersection>291 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-35,291,-29,291</points>
<intersection>-35 0</intersection>
<intersection>-29 1</intersection></hsegment></shape></wire>
<wire>
<ID>1314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,240.5,-50,265.5</points>
<intersection>240.5 1</intersection>
<intersection>265.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,240.5,-45.5,240.5</points>
<connection>
<GID>1411</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1413</GID>
<name>IN_1</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-50,265.5,-44.5,265.5</points>
<intersection>-50 0</intersection>
<intersection>-44.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-44.5,257,-44.5,265.5</points>
<connection>
<GID>1417</GID>
<name>IN_0</name></connection>
<intersection>265.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>1315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,242.5,-63.5,258.5</points>
<intersection>242.5 3</intersection>
<intersection>258.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-79,258.5,-62,258.5</points>
<connection>
<GID>1409</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 0</intersection>
<intersection>-62 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-63.5,242.5,-45.5,242.5</points>
<connection>
<GID>1413</GID>
<name>IN_0</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-62,258,-62,258.5</points>
<connection>
<GID>1415</GID>
<name>IN_0</name></connection>
<intersection>258.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,257,-46.5,258</points>
<connection>
<GID>1417</GID>
<name>IN_1</name></connection>
<intersection>258 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,258,-46.5,258</points>
<connection>
<GID>1415</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45.5,250.5,-40,250.5</points>
<intersection>-45.5 5</intersection>
<intersection>-40 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-40,250.5,-40,255</points>
<intersection>250.5 1</intersection>
<intersection>255 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-45.5,250.5,-45.5,251</points>
<connection>
<GID>1417</GID>
<name>OUT</name></connection>
<intersection>250.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-40,255,-36.5,255</points>
<connection>
<GID>1585</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></hsegment></shape></wire>
<wire>
<ID>1318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,255,-26,271.5</points>
<intersection>255 1</intersection>
<intersection>271.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30.5,255,-26,255</points>
<connection>
<GID>1585</GID>
<name>OUT_0</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26,271.5,43.5,271.5</points>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection>
<intersection>-26 0</intersection></hsegment></shape></wire>
<wire>
<ID>1319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30.5,252,42.5,252</points>
<connection>
<GID>1585</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>1567</GID>
<name>IN_1</name></connection>
<intersection>-5.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-5.5,147.5,-5.5,252</points>
<intersection>147.5 8</intersection>
<intersection>252 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-5.5,147.5,39.5,147.5</points>
<connection>
<GID>1429</GID>
<name>IN_3</name></connection>
<intersection>-5.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39.5,437,603.5,437</points>
<intersection>-39.5 15</intersection>
<intersection>-32 16</intersection>
<intersection>239.5 25</intersection>
<intersection>603.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>603.5,48.5,603.5,437</points>
<intersection>48.5 3</intersection>
<intersection>437 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>446.5,48.5,603.5,48.5</points>
<intersection>446.5 14</intersection>
<intersection>462.5 13</intersection>
<intersection>476 12</intersection>
<intersection>491 11</intersection>
<intersection>501.5 10</intersection>
<intersection>514.5 9</intersection>
<intersection>603.5 2</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>514.5,48.5,514.5,60</points>
<connection>
<GID>1441</GID>
<name>clock</name></connection>
<intersection>48.5 3</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>501.5,48.5,501.5,60</points>
<connection>
<GID>1435</GID>
<name>clock</name></connection>
<intersection>48.5 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>491,48.5,491,60</points>
<connection>
<GID>1430</GID>
<name>clock</name></connection>
<intersection>48.5 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>476,48.5,476,60</points>
<connection>
<GID>1423</GID>
<name>clock</name></connection>
<intersection>48.5 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>462.5,48.5,462.5,60</points>
<connection>
<GID>1414</GID>
<name>clock</name></connection>
<intersection>48.5 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>446.5,48.5,446.5,60.5</points>
<connection>
<GID>1566</GID>
<name>clock</name></connection>
<intersection>48.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-39.5,437,-39.5,447.5</points>
<connection>
<GID>1492</GID>
<name>CLK</name></connection>
<intersection>437 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-32,437,-32,447.5</points>
<connection>
<GID>1462</GID>
<name>IN_1</name></connection>
<intersection>437 1</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>239.5,386,239.5,437</points>
<intersection>386 26</intersection>
<intersection>437 1</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>227,386,239.5,386</points>
<connection>
<GID>1449</GID>
<name>clock</name></connection>
<intersection>239.5 25</intersection></hsegment></shape></wire>
<wire>
<ID>1322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,396.5,-15,401</points>
<intersection>396.5 1</intersection>
<intersection>401 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18.5,396.5,-15,396.5</points>
<connection>
<GID>1467</GID>
<name>IN_1</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,401,-11.5,401</points>
<connection>
<GID>1466</GID>
<name>OUT</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>1324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-24.5,384,205.5,384</points>
<connection>
<GID>1493</GID>
<name>clear</name></connection>
<connection>
<GID>1481</GID>
<name>clear</name></connection>
<connection>
<GID>1483</GID>
<name>clear</name></connection>
<connection>
<GID>1485</GID>
<name>clear</name></connection>
<connection>
<GID>1491</GID>
<name>clear</name></connection>
<connection>
<GID>1460</GID>
<name>OUT</name></connection>
<intersection>-24.5 6</intersection>
<intersection>112 4</intersection>
<intersection>157.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>157.5,383.5,157.5,384</points>
<connection>
<GID>1488</GID>
<name>clear</name></connection>
<intersection>384 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>112,348,112,384</points>
<intersection>348 5</intersection>
<intersection>384 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>112,348,203,348</points>
<intersection>112 4</intersection>
<intersection>121 13</intersection>
<intersection>137.5 12</intersection>
<intersection>152 11</intersection>
<intersection>169 10</intersection>
<intersection>185 9</intersection>
<intersection>203 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-24.5,384,-24.5,404</points>
<intersection>384 1</intersection>
<intersection>404 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-25,404,-24.5,404</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<intersection>-24.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>203,348,203,349</points>
<connection>
<GID>1511</GID>
<name>clear</name></connection>
<intersection>348 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>185,348,185,349</points>
<connection>
<GID>1510</GID>
<name>clear</name></connection>
<intersection>348 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>169,348,169,349</points>
<connection>
<GID>1509</GID>
<name>clear</name></connection>
<intersection>348 5</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>152,348,152,349</points>
<connection>
<GID>1507</GID>
<name>clear</name></connection>
<intersection>348 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>137.5,348,137.5,349</points>
<connection>
<GID>1506</GID>
<name>clear</name></connection>
<intersection>348 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>121,348,121,349</points>
<connection>
<GID>1504</GID>
<name>clear</name></connection>
<intersection>348 5</intersection></vsegment></shape></wire>
<wire>
<ID>1325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18.5,394.5,21.5,394.5</points>
<connection>
<GID>1467</GID>
<name>IN_0</name></connection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,392.5,21.5,394.5</points>
<connection>
<GID>1464</GID>
<name>OUT</name></connection>
<intersection>394.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,405,-37,409</points>
<intersection>405 2</intersection>
<intersection>409 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43.5,409,-37,409</points>
<connection>
<GID>1473</GID>
<name>IN_1</name></connection>
<intersection>-37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37,405,-31,405</points>
<connection>
<GID>1470</GID>
<name>OUT</name></connection>
<intersection>-37 0</intersection></hsegment></shape></wire>
<wire>
<ID>1328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,457,29,457</points>
<connection>
<GID>1471</GID>
<name>clear</name></connection>
<connection>
<GID>1469</GID>
<name>clear</name></connection>
<connection>
<GID>1468</GID>
<name>clear</name></connection>
<intersection>-16.5 13</intersection>
<intersection>29 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29,456,29,457</points>
<connection>
<GID>1474</GID>
<name>clear</name></connection>
<intersection>456 5</intersection>
<intersection>457 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>29,456,110.5,456</points>
<connection>
<GID>1477</GID>
<name>clear</name></connection>
<connection>
<GID>1476</GID>
<name>clear</name></connection>
<intersection>29 4</intersection>
<intersection>91.5 30</intersection>
<intersection>110.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>110.5,449,110.5,456</points>
<connection>
<GID>1513</GID>
<name>IN_0</name></connection>
<intersection>456 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-16.5,422,-16.5,457</points>
<intersection>422 14</intersection>
<intersection>457 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-16.5,422,74.5,422</points>
<connection>
<GID>1519</GID>
<name>clear</name></connection>
<connection>
<GID>1518</GID>
<name>clear</name></connection>
<connection>
<GID>1517</GID>
<name>clear</name></connection>
<connection>
<GID>1516</GID>
<name>clear</name></connection>
<connection>
<GID>1515</GID>
<name>clear</name></connection>
<connection>
<GID>1514</GID>
<name>clear</name></connection>
<intersection>-16.5 13</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>91.5,456,91.5,463</points>
<connection>
<GID>1478</GID>
<name>OUT</name></connection>
<intersection>456 5</intersection></vsegment></shape></wire>
<wire>
<ID>1329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,475.5,112.5,475.5</points>
<intersection>79.5 3</intersection>
<intersection>112.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>79.5,471.5,79.5,475.5</points>
<intersection>471.5 5</intersection>
<intersection>475.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>112.5,473,112.5,475.5</points>
<connection>
<GID>1456</GID>
<name>IN_1</name></connection>
<intersection>475.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>78.5,471.5,79.5,471.5</points>
<connection>
<GID>1508</GID>
<name>OUT</name></connection>
<intersection>79.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,398.5,210.5,401</points>
<intersection>398.5 2</intersection>
<intersection>401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,401,214.5,401</points>
<connection>
<GID>1461</GID>
<name>IN_0</name></connection>
<intersection>210.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,398.5,210.5,398.5</points>
<connection>
<GID>1503</GID>
<name>OUT</name></connection>
<intersection>210.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,395.5,-24.5,395.5</points>
<connection>
<GID>1482</GID>
<name>IN_0</name></connection>
<connection>
<GID>1467</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,396.5,-42,407</points>
<connection>
<GID>1482</GID>
<name>OUT</name></connection>
<intersection>407 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43.5,407,-42,407</points>
<connection>
<GID>1473</GID>
<name>IN_0</name></connection>
<intersection>-42 0</intersection></hsegment></shape></wire>
<wire>
<ID>1334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-57.5,408,-49.5,408</points>
<connection>
<GID>1487</GID>
<name>N_in1</name></connection>
<connection>
<GID>1473</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,464,102,472</points>
<intersection>464 1</intersection>
<intersection>472 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,464,102,464</points>
<connection>
<GID>1478</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,472,106.5,472</points>
<connection>
<GID>1456</GID>
<name>OUT</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>1336</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-36,379.5,211.5,379.5</points>
<connection>
<GID>1465</GID>
<name>OUT_0</name></connection>
<intersection>97.5 15</intersection>
<intersection>211.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>211.5,379.5,211.5,383</points>
<connection>
<GID>1460</GID>
<name>IN_0</name></connection>
<intersection>379.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>97.5,379.5,97.5,462</points>
<connection>
<GID>1478</GID>
<name>IN_0</name></connection>
<intersection>379.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>1337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,459,8.5,471.5</points>
<intersection>459 4</intersection>
<intersection>463 2</intersection>
<intersection>471.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,471.5,18,471.5</points>
<connection>
<GID>1495</GID>
<name>OUT</name></connection>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,463,10,463</points>
<connection>
<GID>1471</GID>
<name>J</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8.5,459,10,459</points>
<connection>
<GID>1471</GID>
<name>K</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,458.5,25,470.5</points>
<intersection>458.5 4</intersection>
<intersection>462.5 2</intersection>
<intersection>470.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,470.5,33,470.5</points>
<connection>
<GID>1499</GID>
<name>OUT</name></connection>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,462.5,26,462.5</points>
<connection>
<GID>1474</GID>
<name>J</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>25,458.5,26,458.5</points>
<connection>
<GID>1474</GID>
<name>K</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>1339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,458,40.5,469.5</points>
<intersection>458 4</intersection>
<intersection>462 2</intersection>
<intersection>469.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,469.5,50.5,469.5</points>
<connection>
<GID>1502</GID>
<name>OUT</name></connection>
<connection>
<GID>1505</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,462,42,462</points>
<connection>
<GID>1476</GID>
<name>J</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40.5,458,42,458</points>
<connection>
<GID>1476</GID>
<name>K</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,458,57.5,468.5</points>
<intersection>458 4</intersection>
<intersection>462 2</intersection>
<intersection>468.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,468.5,57.5,468.5</points>
<connection>
<GID>1505</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,462,59,462</points>
<connection>
<GID>1477</GID>
<name>J</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>57.5,458,59,458</points>
<connection>
<GID>1477</GID>
<name>K</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,463,-6,463</points>
<connection>
<GID>1468</GID>
<name>Q</name></connection>
<connection>
<GID>1469</GID>
<name>J</name></connection>
<intersection>-12.5 3</intersection>
<intersection>-10 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-12.5,428,-12.5,463</points>
<intersection>428 10</intersection>
<intersection>443.5 4</intersection>
<intersection>459 9</intersection>
<intersection>463 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12.5,443.5,74.5,443.5</points>
<connection>
<GID>1484</GID>
<name>IN_0</name></connection>
<intersection>-12.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-10,463,-10,472.5</points>
<intersection>463 1</intersection>
<intersection>472.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-10,472.5,1,472.5</points>
<connection>
<GID>1495</GID>
<name>IN_0</name></connection>
<intersection>-10 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-12.5,459,-6,459</points>
<connection>
<GID>1469</GID>
<name>K</name></connection>
<intersection>-12.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-12.5,428,-10.5,428</points>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>-12.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25.5,453.5,71.5,453.5</points>
<intersection>-25.5 3</intersection>
<intersection>-10 4</intersection>
<intersection>6 32</intersection>
<intersection>7 5</intersection>
<intersection>20.5 31</intersection>
<intersection>23 16</intersection>
<intersection>37.5 30</intersection>
<intersection>39.5 15</intersection>
<intersection>53.5 29</intersection>
<intersection>54.5 18</intersection>
<intersection>71.5 28</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-25.5,425,-25.5,461</points>
<intersection>425 33</intersection>
<intersection>448.5 39</intersection>
<intersection>453.5 1</intersection>
<intersection>461 13</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-10,453.5,-10,461</points>
<intersection>453.5 1</intersection>
<intersection>461 14</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>7,453.5,7,461</points>
<intersection>453.5 1</intersection>
<intersection>461 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>7,461,10,461</points>
<connection>
<GID>1471</GID>
<name>clock</name></connection>
<intersection>7 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-25.5,461,-19.5,461</points>
<connection>
<GID>1468</GID>
<name>clock</name></connection>
<intersection>-25.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-10,461,-6,461</points>
<connection>
<GID>1469</GID>
<name>clock</name></connection>
<intersection>-10 4</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>39.5,453.5,39.5,460</points>
<intersection>453.5 1</intersection>
<intersection>460 21</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>23,453.5,23,460.5</points>
<intersection>453.5 1</intersection>
<intersection>460.5 19</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>54.5,453.5,54.5,460</points>
<intersection>453.5 1</intersection>
<intersection>460 20</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>23,460.5,26,460.5</points>
<connection>
<GID>1474</GID>
<name>clock</name></connection>
<intersection>23 16</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>54.5,460,59,460</points>
<connection>
<GID>1477</GID>
<name>clock</name></connection>
<intersection>54.5 18</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>39.5,460,42,460</points>
<connection>
<GID>1476</GID>
<name>clock</name></connection>
<intersection>39.5 15</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>71.5,425,71.5,453.5</points>
<connection>
<GID>1519</GID>
<name>clock</name></connection>
<intersection>453.5 1</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>53.5,425,53.5,453.5</points>
<connection>
<GID>1518</GID>
<name>clock</name></connection>
<intersection>453.5 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>37.5,425,37.5,453.5</points>
<connection>
<GID>1517</GID>
<name>clock</name></connection>
<intersection>453.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>20.5,425,20.5,453.5</points>
<connection>
<GID>1516</GID>
<name>clock</name></connection>
<intersection>453.5 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>6,425,6,453.5</points>
<connection>
<GID>1515</GID>
<name>clock</name></connection>
<intersection>453.5 1</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-25.5,425,-10.5,425</points>
<connection>
<GID>1514</GID>
<name>clock</name></connection>
<intersection>-25.5 3</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-26,448.5,-25.5,448.5</points>
<connection>
<GID>1462</GID>
<name>OUT</name></connection>
<intersection>-25.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,428,1,470.5</points>
<connection>
<GID>1495</GID>
<name>IN_1</name></connection>
<intersection>428 8</intersection>
<intersection>444.5 1</intersection>
<intersection>463 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,444.5,74.5,444.5</points>
<connection>
<GID>1484</GID>
<name>IN_1</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>0,463,1,463</points>
<connection>
<GID>1469</GID>
<name>Q</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>1,428,6,428</points>
<connection>
<GID>1515</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>1344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,446.5,74.5,446.5</points>
<connection>
<GID>1484</GID>
<name>IN_3</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,428,33,472.5</points>
<connection>
<GID>1502</GID>
<name>IN_1</name></connection>
<intersection>428 9</intersection>
<intersection>446.5 1</intersection>
<intersection>462.5 4</intersection>
<intersection>472.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32,462.5,33,462.5</points>
<connection>
<GID>1474</GID>
<name>Q</name></connection>
<intersection>33 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>33,472.5,72.5,472.5</points>
<connection>
<GID>1508</GID>
<name>IN_1</name></connection>
<intersection>33 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>33,428,37.5,428</points>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>33 3</intersection></hsegment></shape></wire>
<wire>
<ID>1345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,428,17,474.5</points>
<intersection>428 9</intersection>
<intersection>445.5 4</intersection>
<intersection>463 3</intersection>
<intersection>469.5 2</intersection>
<intersection>474.5 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17,469.5,18,469.5</points>
<connection>
<GID>1499</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>16,463,17,463</points>
<connection>
<GID>1471</GID>
<name>Q</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>17,445.5,74.5,445.5</points>
<connection>
<GID>1484</GID>
<name>IN_2</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>17,474.5,72.5,474.5</points>
<connection>
<GID>1508</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>17,428,20.5,428</points>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>1346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,428,49,470.5</points>
<intersection>428 8</intersection>
<intersection>447.5 3</intersection>
<intersection>462 1</intersection>
<intersection>470.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,462,49,462</points>
<connection>
<GID>1476</GID>
<name>Q</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,470.5,72.5,470.5</points>
<connection>
<GID>1508</GID>
<name>IN_2</name></connection>
<intersection>49 0</intersection>
<intersection>50.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>49,447.5,74.5,447.5</points>
<connection>
<GID>1484</GID>
<name>IN_4</name></connection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>50.5,467.5,50.5,470.5</points>
<connection>
<GID>1505</GID>
<name>IN_1</name></connection>
<intersection>470.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>49,428,53.5,428</points>
<connection>
<GID>1518</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>1347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,428,67,468.5</points>
<intersection>428 5</intersection>
<intersection>448.5 2</intersection>
<intersection>462 1</intersection>
<intersection>468.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,462,67,462</points>
<connection>
<GID>1477</GID>
<name>Q</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67,448.5,74.5,448.5</points>
<connection>
<GID>1484</GID>
<name>IN_5</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>67,468.5,72.5,468.5</points>
<connection>
<GID>1508</GID>
<name>IN_3</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>67,428,71.5,428</points>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>1348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3,413.5,89.5,413.5</points>
<connection>
<GID>1520</GID>
<name>IN_0</name></connection>
<intersection>-3 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-3,404,-3,428</points>
<intersection>404 8</intersection>
<intersection>413.5 1</intersection>
<intersection>428 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,428,-3,428</points>
<connection>
<GID>1514</GID>
<name>OUT_0</name></connection>
<intersection>-3 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-4.5,404,-3,404</points>
<connection>
<GID>1466</GID>
<name>IN_3</name></connection>
<intersection>-3 3</intersection></hsegment></shape></wire>
<wire>
<ID>1349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,414.5,89.5,414.5</points>
<connection>
<GID>1520</GID>
<name>IN_1</name></connection>
<intersection>13.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,402,13.5,428</points>
<intersection>402 8</intersection>
<intersection>414.5 1</intersection>
<intersection>428 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>12,428,13.5,428</points>
<connection>
<GID>1515</GID>
<name>OUT_0</name></connection>
<intersection>13.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-4.5,402,13.5,402</points>
<connection>
<GID>1466</GID>
<name>IN_2</name></connection>
<intersection>13.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,415.5,89.5,415.5</points>
<connection>
<GID>1520</GID>
<name>IN_2</name></connection>
<intersection>27.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,400,27.5,428</points>
<intersection>400 8</intersection>
<intersection>415.5 1</intersection>
<intersection>428 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26.5,428,27.5,428</points>
<connection>
<GID>1516</GID>
<name>OUT_0</name></connection>
<intersection>27.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-4.5,400,27.5,400</points>
<connection>
<GID>1466</GID>
<name>IN_1</name></connection>
<intersection>27.5 3</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>-83.0729,339.455,1140.93,-265.545</PageViewport></page 6>
<page 7>
<PageViewport>-83.0729,339.455,1140.93,-265.545</PageViewport></page 7>
<page 8>
<PageViewport>-83.0729,339.455,1140.93,-265.545</PageViewport></page 8>
<page 9>
<PageViewport>-83.0729,339.455,1140.93,-265.545</PageViewport></page 9></circuit>